magic
tech gf180mcuC
magscale 1 10
timestamp 1670141033
<< obsm1 >>
rect 1344 1710 579134 579570
<< metal2 >>
rect 9296 582153 9408 582953
rect 25312 582153 25424 582953
rect 41328 582153 41440 582953
rect 57344 582153 57456 582953
rect 73360 582153 73472 582953
rect 89376 582153 89488 582953
rect 105392 582153 105504 582953
rect 121408 582153 121520 582953
rect 137424 582153 137536 582953
rect 153440 582153 153552 582953
rect 169456 582153 169568 582953
rect 185472 582153 185584 582953
rect 201488 582153 201600 582953
rect 217504 582153 217616 582953
rect 233520 582153 233632 582953
rect 249536 582153 249648 582953
rect 265552 582153 265664 582953
rect 281568 582153 281680 582953
rect 297584 582153 297696 582953
rect 313600 582153 313712 582953
rect 329616 582153 329728 582953
rect 345632 582153 345744 582953
rect 361648 582153 361760 582953
rect 377664 582153 377776 582953
rect 393680 582153 393792 582953
rect 409696 582153 409808 582953
rect 425712 582153 425824 582953
rect 441728 582153 441840 582953
rect 457744 582153 457856 582953
rect 473760 582153 473872 582953
rect 489776 582153 489888 582953
rect 505792 582153 505904 582953
rect 521808 582153 521920 582953
rect 537824 582153 537936 582953
rect 553840 582153 553952 582953
rect 569856 582153 569968 582953
rect 3024 0 3136 800
rect 4928 0 5040 800
rect 6832 0 6944 800
rect 8736 0 8848 800
rect 10640 0 10752 800
rect 12544 0 12656 800
rect 14448 0 14560 800
rect 16352 0 16464 800
rect 18256 0 18368 800
rect 20160 0 20272 800
rect 22064 0 22176 800
rect 23968 0 24080 800
rect 25872 0 25984 800
rect 27776 0 27888 800
rect 29680 0 29792 800
rect 31584 0 31696 800
rect 33488 0 33600 800
rect 35392 0 35504 800
rect 37296 0 37408 800
rect 39200 0 39312 800
rect 41104 0 41216 800
rect 43008 0 43120 800
rect 44912 0 45024 800
rect 46816 0 46928 800
rect 48720 0 48832 800
rect 50624 0 50736 800
rect 52528 0 52640 800
rect 54432 0 54544 800
rect 56336 0 56448 800
rect 58240 0 58352 800
rect 60144 0 60256 800
rect 62048 0 62160 800
rect 63952 0 64064 800
rect 65856 0 65968 800
rect 67760 0 67872 800
rect 69664 0 69776 800
rect 71568 0 71680 800
rect 73472 0 73584 800
rect 75376 0 75488 800
rect 77280 0 77392 800
rect 79184 0 79296 800
rect 81088 0 81200 800
rect 82992 0 83104 800
rect 84896 0 85008 800
rect 86800 0 86912 800
rect 88704 0 88816 800
rect 90608 0 90720 800
rect 92512 0 92624 800
rect 94416 0 94528 800
rect 96320 0 96432 800
rect 98224 0 98336 800
rect 100128 0 100240 800
rect 102032 0 102144 800
rect 103936 0 104048 800
rect 105840 0 105952 800
rect 107744 0 107856 800
rect 109648 0 109760 800
rect 111552 0 111664 800
rect 113456 0 113568 800
rect 115360 0 115472 800
rect 117264 0 117376 800
rect 119168 0 119280 800
rect 121072 0 121184 800
rect 122976 0 123088 800
rect 124880 0 124992 800
rect 126784 0 126896 800
rect 128688 0 128800 800
rect 130592 0 130704 800
rect 132496 0 132608 800
rect 134400 0 134512 800
rect 136304 0 136416 800
rect 138208 0 138320 800
rect 140112 0 140224 800
rect 142016 0 142128 800
rect 143920 0 144032 800
rect 145824 0 145936 800
rect 147728 0 147840 800
rect 149632 0 149744 800
rect 151536 0 151648 800
rect 153440 0 153552 800
rect 155344 0 155456 800
rect 157248 0 157360 800
rect 159152 0 159264 800
rect 161056 0 161168 800
rect 162960 0 163072 800
rect 164864 0 164976 800
rect 166768 0 166880 800
rect 168672 0 168784 800
rect 170576 0 170688 800
rect 172480 0 172592 800
rect 174384 0 174496 800
rect 176288 0 176400 800
rect 178192 0 178304 800
rect 180096 0 180208 800
rect 182000 0 182112 800
rect 183904 0 184016 800
rect 185808 0 185920 800
rect 187712 0 187824 800
rect 189616 0 189728 800
rect 191520 0 191632 800
rect 193424 0 193536 800
rect 195328 0 195440 800
rect 197232 0 197344 800
rect 199136 0 199248 800
rect 201040 0 201152 800
rect 202944 0 203056 800
rect 204848 0 204960 800
rect 206752 0 206864 800
rect 208656 0 208768 800
rect 210560 0 210672 800
rect 212464 0 212576 800
rect 214368 0 214480 800
rect 216272 0 216384 800
rect 218176 0 218288 800
rect 220080 0 220192 800
rect 221984 0 222096 800
rect 223888 0 224000 800
rect 225792 0 225904 800
rect 227696 0 227808 800
rect 229600 0 229712 800
rect 231504 0 231616 800
rect 233408 0 233520 800
rect 235312 0 235424 800
rect 237216 0 237328 800
rect 239120 0 239232 800
rect 241024 0 241136 800
rect 242928 0 243040 800
rect 244832 0 244944 800
rect 246736 0 246848 800
rect 248640 0 248752 800
rect 250544 0 250656 800
rect 252448 0 252560 800
rect 254352 0 254464 800
rect 256256 0 256368 800
rect 258160 0 258272 800
rect 260064 0 260176 800
rect 261968 0 262080 800
rect 263872 0 263984 800
rect 265776 0 265888 800
rect 267680 0 267792 800
rect 269584 0 269696 800
rect 271488 0 271600 800
rect 273392 0 273504 800
rect 275296 0 275408 800
rect 277200 0 277312 800
rect 279104 0 279216 800
rect 281008 0 281120 800
rect 282912 0 283024 800
rect 284816 0 284928 800
rect 286720 0 286832 800
rect 288624 0 288736 800
rect 290528 0 290640 800
rect 292432 0 292544 800
rect 294336 0 294448 800
rect 296240 0 296352 800
rect 298144 0 298256 800
rect 300048 0 300160 800
rect 301952 0 302064 800
rect 303856 0 303968 800
rect 305760 0 305872 800
rect 307664 0 307776 800
rect 309568 0 309680 800
rect 311472 0 311584 800
rect 313376 0 313488 800
rect 315280 0 315392 800
rect 317184 0 317296 800
rect 319088 0 319200 800
rect 320992 0 321104 800
rect 322896 0 323008 800
rect 324800 0 324912 800
rect 326704 0 326816 800
rect 328608 0 328720 800
rect 330512 0 330624 800
rect 332416 0 332528 800
rect 334320 0 334432 800
rect 336224 0 336336 800
rect 338128 0 338240 800
rect 340032 0 340144 800
rect 341936 0 342048 800
rect 343840 0 343952 800
rect 345744 0 345856 800
rect 347648 0 347760 800
rect 349552 0 349664 800
rect 351456 0 351568 800
rect 353360 0 353472 800
rect 355264 0 355376 800
rect 357168 0 357280 800
rect 359072 0 359184 800
rect 360976 0 361088 800
rect 362880 0 362992 800
rect 364784 0 364896 800
rect 366688 0 366800 800
rect 368592 0 368704 800
rect 370496 0 370608 800
rect 372400 0 372512 800
rect 374304 0 374416 800
rect 376208 0 376320 800
rect 378112 0 378224 800
rect 380016 0 380128 800
rect 381920 0 382032 800
rect 383824 0 383936 800
rect 385728 0 385840 800
rect 387632 0 387744 800
rect 389536 0 389648 800
rect 391440 0 391552 800
rect 393344 0 393456 800
rect 395248 0 395360 800
rect 397152 0 397264 800
rect 399056 0 399168 800
rect 400960 0 401072 800
rect 402864 0 402976 800
rect 404768 0 404880 800
rect 406672 0 406784 800
rect 408576 0 408688 800
rect 410480 0 410592 800
rect 412384 0 412496 800
rect 414288 0 414400 800
rect 416192 0 416304 800
rect 418096 0 418208 800
rect 420000 0 420112 800
rect 421904 0 422016 800
rect 423808 0 423920 800
rect 425712 0 425824 800
rect 427616 0 427728 800
rect 429520 0 429632 800
rect 431424 0 431536 800
rect 433328 0 433440 800
rect 435232 0 435344 800
rect 437136 0 437248 800
rect 439040 0 439152 800
rect 440944 0 441056 800
rect 442848 0 442960 800
rect 444752 0 444864 800
rect 446656 0 446768 800
rect 448560 0 448672 800
rect 450464 0 450576 800
rect 452368 0 452480 800
rect 454272 0 454384 800
rect 456176 0 456288 800
rect 458080 0 458192 800
rect 459984 0 460096 800
rect 461888 0 462000 800
rect 463792 0 463904 800
rect 465696 0 465808 800
rect 467600 0 467712 800
rect 469504 0 469616 800
rect 471408 0 471520 800
rect 473312 0 473424 800
rect 475216 0 475328 800
rect 477120 0 477232 800
rect 479024 0 479136 800
rect 480928 0 481040 800
rect 482832 0 482944 800
rect 484736 0 484848 800
rect 486640 0 486752 800
rect 488544 0 488656 800
rect 490448 0 490560 800
rect 492352 0 492464 800
rect 494256 0 494368 800
rect 496160 0 496272 800
rect 498064 0 498176 800
rect 499968 0 500080 800
rect 501872 0 501984 800
rect 503776 0 503888 800
rect 505680 0 505792 800
rect 507584 0 507696 800
rect 509488 0 509600 800
rect 511392 0 511504 800
rect 513296 0 513408 800
rect 515200 0 515312 800
rect 517104 0 517216 800
rect 519008 0 519120 800
rect 520912 0 521024 800
rect 522816 0 522928 800
rect 524720 0 524832 800
rect 526624 0 526736 800
rect 528528 0 528640 800
rect 530432 0 530544 800
rect 532336 0 532448 800
rect 534240 0 534352 800
rect 536144 0 536256 800
rect 538048 0 538160 800
rect 539952 0 540064 800
rect 541856 0 541968 800
rect 543760 0 543872 800
rect 545664 0 545776 800
rect 547568 0 547680 800
rect 549472 0 549584 800
rect 551376 0 551488 800
rect 553280 0 553392 800
rect 555184 0 555296 800
rect 557088 0 557200 800
rect 558992 0 559104 800
rect 560896 0 561008 800
rect 562800 0 562912 800
rect 564704 0 564816 800
rect 566608 0 566720 800
rect 568512 0 568624 800
rect 570416 0 570528 800
rect 572320 0 572432 800
rect 574224 0 574336 800
rect 576128 0 576240 800
<< obsm2 >>
rect 812 582093 9236 582153
rect 9468 582093 25252 582153
rect 25484 582093 41268 582153
rect 41500 582093 57284 582153
rect 57516 582093 73300 582153
rect 73532 582093 89316 582153
rect 89548 582093 105332 582153
rect 105564 582093 121348 582153
rect 121580 582093 137364 582153
rect 137596 582093 153380 582153
rect 153612 582093 169396 582153
rect 169628 582093 185412 582153
rect 185644 582093 201428 582153
rect 201660 582093 217444 582153
rect 217676 582093 233460 582153
rect 233692 582093 249476 582153
rect 249708 582093 265492 582153
rect 265724 582093 281508 582153
rect 281740 582093 297524 582153
rect 297756 582093 313540 582153
rect 313772 582093 329556 582153
rect 329788 582093 345572 582153
rect 345804 582093 361588 582153
rect 361820 582093 377604 582153
rect 377836 582093 393620 582153
rect 393852 582093 409636 582153
rect 409868 582093 425652 582153
rect 425884 582093 441668 582153
rect 441900 582093 457684 582153
rect 457916 582093 473700 582153
rect 473932 582093 489716 582153
rect 489948 582093 505732 582153
rect 505964 582093 521748 582153
rect 521980 582093 537764 582153
rect 537996 582093 553780 582153
rect 554012 582093 569796 582153
rect 570028 582093 579348 582153
rect 812 860 579348 582093
rect 812 354 2964 860
rect 3196 354 4868 860
rect 5100 354 6772 860
rect 7004 354 8676 860
rect 8908 354 10580 860
rect 10812 354 12484 860
rect 12716 354 14388 860
rect 14620 354 16292 860
rect 16524 354 18196 860
rect 18428 354 20100 860
rect 20332 354 22004 860
rect 22236 354 23908 860
rect 24140 354 25812 860
rect 26044 354 27716 860
rect 27948 354 29620 860
rect 29852 354 31524 860
rect 31756 354 33428 860
rect 33660 354 35332 860
rect 35564 354 37236 860
rect 37468 354 39140 860
rect 39372 354 41044 860
rect 41276 354 42948 860
rect 43180 354 44852 860
rect 45084 354 46756 860
rect 46988 354 48660 860
rect 48892 354 50564 860
rect 50796 354 52468 860
rect 52700 354 54372 860
rect 54604 354 56276 860
rect 56508 354 58180 860
rect 58412 354 60084 860
rect 60316 354 61988 860
rect 62220 354 63892 860
rect 64124 354 65796 860
rect 66028 354 67700 860
rect 67932 354 69604 860
rect 69836 354 71508 860
rect 71740 354 73412 860
rect 73644 354 75316 860
rect 75548 354 77220 860
rect 77452 354 79124 860
rect 79356 354 81028 860
rect 81260 354 82932 860
rect 83164 354 84836 860
rect 85068 354 86740 860
rect 86972 354 88644 860
rect 88876 354 90548 860
rect 90780 354 92452 860
rect 92684 354 94356 860
rect 94588 354 96260 860
rect 96492 354 98164 860
rect 98396 354 100068 860
rect 100300 354 101972 860
rect 102204 354 103876 860
rect 104108 354 105780 860
rect 106012 354 107684 860
rect 107916 354 109588 860
rect 109820 354 111492 860
rect 111724 354 113396 860
rect 113628 354 115300 860
rect 115532 354 117204 860
rect 117436 354 119108 860
rect 119340 354 121012 860
rect 121244 354 122916 860
rect 123148 354 124820 860
rect 125052 354 126724 860
rect 126956 354 128628 860
rect 128860 354 130532 860
rect 130764 354 132436 860
rect 132668 354 134340 860
rect 134572 354 136244 860
rect 136476 354 138148 860
rect 138380 354 140052 860
rect 140284 354 141956 860
rect 142188 354 143860 860
rect 144092 354 145764 860
rect 145996 354 147668 860
rect 147900 354 149572 860
rect 149804 354 151476 860
rect 151708 354 153380 860
rect 153612 354 155284 860
rect 155516 354 157188 860
rect 157420 354 159092 860
rect 159324 354 160996 860
rect 161228 354 162900 860
rect 163132 354 164804 860
rect 165036 354 166708 860
rect 166940 354 168612 860
rect 168844 354 170516 860
rect 170748 354 172420 860
rect 172652 354 174324 860
rect 174556 354 176228 860
rect 176460 354 178132 860
rect 178364 354 180036 860
rect 180268 354 181940 860
rect 182172 354 183844 860
rect 184076 354 185748 860
rect 185980 354 187652 860
rect 187884 354 189556 860
rect 189788 354 191460 860
rect 191692 354 193364 860
rect 193596 354 195268 860
rect 195500 354 197172 860
rect 197404 354 199076 860
rect 199308 354 200980 860
rect 201212 354 202884 860
rect 203116 354 204788 860
rect 205020 354 206692 860
rect 206924 354 208596 860
rect 208828 354 210500 860
rect 210732 354 212404 860
rect 212636 354 214308 860
rect 214540 354 216212 860
rect 216444 354 218116 860
rect 218348 354 220020 860
rect 220252 354 221924 860
rect 222156 354 223828 860
rect 224060 354 225732 860
rect 225964 354 227636 860
rect 227868 354 229540 860
rect 229772 354 231444 860
rect 231676 354 233348 860
rect 233580 354 235252 860
rect 235484 354 237156 860
rect 237388 354 239060 860
rect 239292 354 240964 860
rect 241196 354 242868 860
rect 243100 354 244772 860
rect 245004 354 246676 860
rect 246908 354 248580 860
rect 248812 354 250484 860
rect 250716 354 252388 860
rect 252620 354 254292 860
rect 254524 354 256196 860
rect 256428 354 258100 860
rect 258332 354 260004 860
rect 260236 354 261908 860
rect 262140 354 263812 860
rect 264044 354 265716 860
rect 265948 354 267620 860
rect 267852 354 269524 860
rect 269756 354 271428 860
rect 271660 354 273332 860
rect 273564 354 275236 860
rect 275468 354 277140 860
rect 277372 354 279044 860
rect 279276 354 280948 860
rect 281180 354 282852 860
rect 283084 354 284756 860
rect 284988 354 286660 860
rect 286892 354 288564 860
rect 288796 354 290468 860
rect 290700 354 292372 860
rect 292604 354 294276 860
rect 294508 354 296180 860
rect 296412 354 298084 860
rect 298316 354 299988 860
rect 300220 354 301892 860
rect 302124 354 303796 860
rect 304028 354 305700 860
rect 305932 354 307604 860
rect 307836 354 309508 860
rect 309740 354 311412 860
rect 311644 354 313316 860
rect 313548 354 315220 860
rect 315452 354 317124 860
rect 317356 354 319028 860
rect 319260 354 320932 860
rect 321164 354 322836 860
rect 323068 354 324740 860
rect 324972 354 326644 860
rect 326876 354 328548 860
rect 328780 354 330452 860
rect 330684 354 332356 860
rect 332588 354 334260 860
rect 334492 354 336164 860
rect 336396 354 338068 860
rect 338300 354 339972 860
rect 340204 354 341876 860
rect 342108 354 343780 860
rect 344012 354 345684 860
rect 345916 354 347588 860
rect 347820 354 349492 860
rect 349724 354 351396 860
rect 351628 354 353300 860
rect 353532 354 355204 860
rect 355436 354 357108 860
rect 357340 354 359012 860
rect 359244 354 360916 860
rect 361148 354 362820 860
rect 363052 354 364724 860
rect 364956 354 366628 860
rect 366860 354 368532 860
rect 368764 354 370436 860
rect 370668 354 372340 860
rect 372572 354 374244 860
rect 374476 354 376148 860
rect 376380 354 378052 860
rect 378284 354 379956 860
rect 380188 354 381860 860
rect 382092 354 383764 860
rect 383996 354 385668 860
rect 385900 354 387572 860
rect 387804 354 389476 860
rect 389708 354 391380 860
rect 391612 354 393284 860
rect 393516 354 395188 860
rect 395420 354 397092 860
rect 397324 354 398996 860
rect 399228 354 400900 860
rect 401132 354 402804 860
rect 403036 354 404708 860
rect 404940 354 406612 860
rect 406844 354 408516 860
rect 408748 354 410420 860
rect 410652 354 412324 860
rect 412556 354 414228 860
rect 414460 354 416132 860
rect 416364 354 418036 860
rect 418268 354 419940 860
rect 420172 354 421844 860
rect 422076 354 423748 860
rect 423980 354 425652 860
rect 425884 354 427556 860
rect 427788 354 429460 860
rect 429692 354 431364 860
rect 431596 354 433268 860
rect 433500 354 435172 860
rect 435404 354 437076 860
rect 437308 354 438980 860
rect 439212 354 440884 860
rect 441116 354 442788 860
rect 443020 354 444692 860
rect 444924 354 446596 860
rect 446828 354 448500 860
rect 448732 354 450404 860
rect 450636 354 452308 860
rect 452540 354 454212 860
rect 454444 354 456116 860
rect 456348 354 458020 860
rect 458252 354 459924 860
rect 460156 354 461828 860
rect 462060 354 463732 860
rect 463964 354 465636 860
rect 465868 354 467540 860
rect 467772 354 469444 860
rect 469676 354 471348 860
rect 471580 354 473252 860
rect 473484 354 475156 860
rect 475388 354 477060 860
rect 477292 354 478964 860
rect 479196 354 480868 860
rect 481100 354 482772 860
rect 483004 354 484676 860
rect 484908 354 486580 860
rect 486812 354 488484 860
rect 488716 354 490388 860
rect 490620 354 492292 860
rect 492524 354 494196 860
rect 494428 354 496100 860
rect 496332 354 498004 860
rect 498236 354 499908 860
rect 500140 354 501812 860
rect 502044 354 503716 860
rect 503948 354 505620 860
rect 505852 354 507524 860
rect 507756 354 509428 860
rect 509660 354 511332 860
rect 511564 354 513236 860
rect 513468 354 515140 860
rect 515372 354 517044 860
rect 517276 354 518948 860
rect 519180 354 520852 860
rect 521084 354 522756 860
rect 522988 354 524660 860
rect 524892 354 526564 860
rect 526796 354 528468 860
rect 528700 354 530372 860
rect 530604 354 532276 860
rect 532508 354 534180 860
rect 534412 354 536084 860
rect 536316 354 537988 860
rect 538220 354 539892 860
rect 540124 354 541796 860
rect 542028 354 543700 860
rect 543932 354 545604 860
rect 545836 354 547508 860
rect 547740 354 549412 860
rect 549644 354 551316 860
rect 551548 354 553220 860
rect 553452 354 555124 860
rect 555356 354 557028 860
rect 557260 354 558932 860
rect 559164 354 560836 860
rect 561068 354 562740 860
rect 562972 354 564644 860
rect 564876 354 566548 860
rect 566780 354 568452 860
rect 568684 354 570356 860
rect 570588 354 572260 860
rect 572492 354 574164 860
rect 574396 354 576068 860
rect 576300 354 579348 860
<< metal3 >>
rect 578569 576800 579369 576912
rect 0 576352 800 576464
rect 578569 565824 579369 565936
rect 0 565600 800 565712
rect 0 554848 800 554960
rect 578569 554848 579369 554960
rect 0 544096 800 544208
rect 578569 543872 579369 543984
rect 0 533344 800 533456
rect 578569 532896 579369 533008
rect 0 522592 800 522704
rect 578569 521920 579369 522032
rect 0 511840 800 511952
rect 578569 510944 579369 511056
rect 0 501088 800 501200
rect 578569 499968 579369 500080
rect 0 490336 800 490448
rect 578569 488992 579369 489104
rect 0 479584 800 479696
rect 578569 478016 579369 478128
rect 0 468832 800 468944
rect 578569 467040 579369 467152
rect 0 458080 800 458192
rect 578569 456064 579369 456176
rect 0 447328 800 447440
rect 578569 445088 579369 445200
rect 0 436576 800 436688
rect 578569 434112 579369 434224
rect 0 425824 800 425936
rect 578569 423136 579369 423248
rect 0 415072 800 415184
rect 578569 412160 579369 412272
rect 0 404320 800 404432
rect 578569 401184 579369 401296
rect 0 393568 800 393680
rect 578569 390208 579369 390320
rect 0 382816 800 382928
rect 578569 379232 579369 379344
rect 0 372064 800 372176
rect 578569 368256 579369 368368
rect 0 361312 800 361424
rect 578569 357280 579369 357392
rect 0 350560 800 350672
rect 578569 346304 579369 346416
rect 0 339808 800 339920
rect 578569 335328 579369 335440
rect 0 329056 800 329168
rect 578569 324352 579369 324464
rect 0 318304 800 318416
rect 578569 313376 579369 313488
rect 0 307552 800 307664
rect 578569 302400 579369 302512
rect 0 296800 800 296912
rect 578569 291424 579369 291536
rect 0 286048 800 286160
rect 578569 280448 579369 280560
rect 0 275296 800 275408
rect 578569 269472 579369 269584
rect 0 264544 800 264656
rect 578569 258496 579369 258608
rect 0 253792 800 253904
rect 578569 247520 579369 247632
rect 0 243040 800 243152
rect 578569 236544 579369 236656
rect 0 232288 800 232400
rect 578569 225568 579369 225680
rect 0 221536 800 221648
rect 578569 214592 579369 214704
rect 0 210784 800 210896
rect 578569 203616 579369 203728
rect 0 200032 800 200144
rect 578569 192640 579369 192752
rect 0 189280 800 189392
rect 578569 181664 579369 181776
rect 0 178528 800 178640
rect 578569 170688 579369 170800
rect 0 167776 800 167888
rect 578569 159712 579369 159824
rect 0 157024 800 157136
rect 578569 148736 579369 148848
rect 0 146272 800 146384
rect 578569 137760 579369 137872
rect 0 135520 800 135632
rect 578569 126784 579369 126896
rect 0 124768 800 124880
rect 578569 115808 579369 115920
rect 0 114016 800 114128
rect 578569 104832 579369 104944
rect 0 103264 800 103376
rect 578569 93856 579369 93968
rect 0 92512 800 92624
rect 578569 82880 579369 82992
rect 0 81760 800 81872
rect 578569 71904 579369 72016
rect 0 71008 800 71120
rect 578569 60928 579369 61040
rect 0 60256 800 60368
rect 578569 49952 579369 50064
rect 0 49504 800 49616
rect 578569 38976 579369 39088
rect 0 38752 800 38864
rect 0 28000 800 28112
rect 578569 28000 579369 28112
rect 0 17248 800 17360
rect 578569 17024 579369 17136
rect 0 6496 800 6608
rect 578569 6048 579369 6160
<< obsm3 >>
rect 800 576972 579358 581252
rect 800 576740 578509 576972
rect 800 576524 579358 576740
rect 860 576292 579358 576524
rect 800 565996 579358 576292
rect 800 565772 578509 565996
rect 860 565764 578509 565772
rect 860 565540 579358 565764
rect 800 555020 579358 565540
rect 860 554788 578509 555020
rect 800 544268 579358 554788
rect 860 544044 579358 544268
rect 860 544036 578509 544044
rect 800 543812 578509 544036
rect 800 533516 579358 543812
rect 860 533284 579358 533516
rect 800 533068 579358 533284
rect 800 532836 578509 533068
rect 800 522764 579358 532836
rect 860 522532 579358 522764
rect 800 522092 579358 522532
rect 800 521860 578509 522092
rect 800 512012 579358 521860
rect 860 511780 579358 512012
rect 800 511116 579358 511780
rect 800 510884 578509 511116
rect 800 501260 579358 510884
rect 860 501028 579358 501260
rect 800 500140 579358 501028
rect 800 499908 578509 500140
rect 800 490508 579358 499908
rect 860 490276 579358 490508
rect 800 489164 579358 490276
rect 800 488932 578509 489164
rect 800 479756 579358 488932
rect 860 479524 579358 479756
rect 800 478188 579358 479524
rect 800 477956 578509 478188
rect 800 469004 579358 477956
rect 860 468772 579358 469004
rect 800 467212 579358 468772
rect 800 466980 578509 467212
rect 800 458252 579358 466980
rect 860 458020 579358 458252
rect 800 456236 579358 458020
rect 800 456004 578509 456236
rect 800 447500 579358 456004
rect 860 447268 579358 447500
rect 800 445260 579358 447268
rect 800 445028 578509 445260
rect 800 436748 579358 445028
rect 860 436516 579358 436748
rect 800 434284 579358 436516
rect 800 434052 578509 434284
rect 800 425996 579358 434052
rect 860 425764 579358 425996
rect 800 423308 579358 425764
rect 800 423076 578509 423308
rect 800 415244 579358 423076
rect 860 415012 579358 415244
rect 800 412332 579358 415012
rect 800 412100 578509 412332
rect 800 404492 579358 412100
rect 860 404260 579358 404492
rect 800 401356 579358 404260
rect 800 401124 578509 401356
rect 800 393740 579358 401124
rect 860 393508 579358 393740
rect 800 390380 579358 393508
rect 800 390148 578509 390380
rect 800 382988 579358 390148
rect 860 382756 579358 382988
rect 800 379404 579358 382756
rect 800 379172 578509 379404
rect 800 372236 579358 379172
rect 860 372004 579358 372236
rect 800 368428 579358 372004
rect 800 368196 578509 368428
rect 800 361484 579358 368196
rect 860 361252 579358 361484
rect 800 357452 579358 361252
rect 800 357220 578509 357452
rect 800 350732 579358 357220
rect 860 350500 579358 350732
rect 800 346476 579358 350500
rect 800 346244 578509 346476
rect 800 339980 579358 346244
rect 860 339748 579358 339980
rect 800 335500 579358 339748
rect 800 335268 578509 335500
rect 800 329228 579358 335268
rect 860 328996 579358 329228
rect 800 324524 579358 328996
rect 800 324292 578509 324524
rect 800 318476 579358 324292
rect 860 318244 579358 318476
rect 800 313548 579358 318244
rect 800 313316 578509 313548
rect 800 307724 579358 313316
rect 860 307492 579358 307724
rect 800 302572 579358 307492
rect 800 302340 578509 302572
rect 800 296972 579358 302340
rect 860 296740 579358 296972
rect 800 291596 579358 296740
rect 800 291364 578509 291596
rect 800 286220 579358 291364
rect 860 285988 579358 286220
rect 800 280620 579358 285988
rect 800 280388 578509 280620
rect 800 275468 579358 280388
rect 860 275236 579358 275468
rect 800 269644 579358 275236
rect 800 269412 578509 269644
rect 800 264716 579358 269412
rect 860 264484 579358 264716
rect 800 258668 579358 264484
rect 800 258436 578509 258668
rect 800 253964 579358 258436
rect 860 253732 579358 253964
rect 800 247692 579358 253732
rect 800 247460 578509 247692
rect 800 243212 579358 247460
rect 860 242980 579358 243212
rect 800 236716 579358 242980
rect 800 236484 578509 236716
rect 800 232460 579358 236484
rect 860 232228 579358 232460
rect 800 225740 579358 232228
rect 800 225508 578509 225740
rect 800 221708 579358 225508
rect 860 221476 579358 221708
rect 800 214764 579358 221476
rect 800 214532 578509 214764
rect 800 210956 579358 214532
rect 860 210724 579358 210956
rect 800 203788 579358 210724
rect 800 203556 578509 203788
rect 800 200204 579358 203556
rect 860 199972 579358 200204
rect 800 192812 579358 199972
rect 800 192580 578509 192812
rect 800 189452 579358 192580
rect 860 189220 579358 189452
rect 800 181836 579358 189220
rect 800 181604 578509 181836
rect 800 178700 579358 181604
rect 860 178468 579358 178700
rect 800 170860 579358 178468
rect 800 170628 578509 170860
rect 800 167948 579358 170628
rect 860 167716 579358 167948
rect 800 159884 579358 167716
rect 800 159652 578509 159884
rect 800 157196 579358 159652
rect 860 156964 579358 157196
rect 800 148908 579358 156964
rect 800 148676 578509 148908
rect 800 146444 579358 148676
rect 860 146212 579358 146444
rect 800 137932 579358 146212
rect 800 137700 578509 137932
rect 800 135692 579358 137700
rect 860 135460 579358 135692
rect 800 126956 579358 135460
rect 800 126724 578509 126956
rect 800 124940 579358 126724
rect 860 124708 579358 124940
rect 800 115980 579358 124708
rect 800 115748 578509 115980
rect 800 114188 579358 115748
rect 860 113956 579358 114188
rect 800 105004 579358 113956
rect 800 104772 578509 105004
rect 800 103436 579358 104772
rect 860 103204 579358 103436
rect 800 94028 579358 103204
rect 800 93796 578509 94028
rect 800 92684 579358 93796
rect 860 92452 579358 92684
rect 800 83052 579358 92452
rect 800 82820 578509 83052
rect 800 81932 579358 82820
rect 860 81700 579358 81932
rect 800 72076 579358 81700
rect 800 71844 578509 72076
rect 800 71180 579358 71844
rect 860 70948 579358 71180
rect 800 61100 579358 70948
rect 800 60868 578509 61100
rect 800 60428 579358 60868
rect 860 60196 579358 60428
rect 800 50124 579358 60196
rect 800 49892 578509 50124
rect 800 49676 579358 49892
rect 860 49444 579358 49676
rect 800 39148 579358 49444
rect 800 38924 578509 39148
rect 860 38916 578509 38924
rect 860 38692 579358 38916
rect 800 28172 579358 38692
rect 860 27940 578509 28172
rect 800 17420 579358 27940
rect 860 17196 579358 17420
rect 860 17188 578509 17196
rect 800 16964 578509 17188
rect 800 6668 579358 16964
rect 860 6436 579358 6668
rect 800 6220 579358 6436
rect 800 5988 578509 6220
rect 800 364 579358 5988
<< metal4 >>
rect 4448 3076 4768 579436
rect 19808 3076 20128 579436
rect 35168 3076 35488 579436
rect 50528 3076 50848 579436
rect 65888 3076 66208 579436
rect 81248 3076 81568 579436
rect 96608 3076 96928 579436
rect 111968 3076 112288 579436
rect 127328 3076 127648 579436
rect 142688 3076 143008 579436
rect 158048 3076 158368 579436
rect 173408 3076 173728 579436
rect 188768 3076 189088 579436
rect 204128 3076 204448 579436
rect 219488 3076 219808 579436
rect 234848 3076 235168 579436
rect 250208 3076 250528 579436
rect 265568 3076 265888 579436
rect 280928 3076 281248 579436
rect 296288 3076 296608 579436
rect 311648 3076 311968 579436
rect 327008 3076 327328 579436
rect 342368 3076 342688 579436
rect 357728 3076 358048 579436
rect 373088 3076 373408 579436
rect 388448 3076 388768 579436
rect 403808 3076 404128 579436
rect 419168 3076 419488 579436
rect 434528 3076 434848 579436
rect 449888 3076 450208 579436
rect 465248 3076 465568 579436
rect 480608 3076 480928 579436
rect 495968 3076 496288 579436
rect 511328 3076 511648 579436
rect 526688 3076 527008 579436
rect 542048 3076 542368 579436
rect 557408 3076 557728 579436
rect 572768 3076 573088 579436
<< obsm4 >>
rect 2380 579496 579348 581150
rect 2380 3016 4388 579496
rect 4828 3016 19748 579496
rect 20188 3016 35108 579496
rect 35548 3016 50468 579496
rect 50908 3016 65828 579496
rect 66268 3016 81188 579496
rect 81628 3016 96548 579496
rect 96988 3016 111908 579496
rect 112348 3016 127268 579496
rect 127708 3016 142628 579496
rect 143068 3016 157988 579496
rect 158428 3016 173348 579496
rect 173788 3016 188708 579496
rect 189148 3016 204068 579496
rect 204508 3016 219428 579496
rect 219868 3016 234788 579496
rect 235228 3016 250148 579496
rect 250588 3016 265508 579496
rect 265948 3016 280868 579496
rect 281308 3016 296228 579496
rect 296668 3016 311588 579496
rect 312028 3016 326948 579496
rect 327388 3016 342308 579496
rect 342748 3016 357668 579496
rect 358108 3016 373028 579496
rect 373468 3016 388388 579496
rect 388828 3016 403748 579496
rect 404188 3016 419108 579496
rect 419548 3016 434468 579496
rect 434908 3016 449828 579496
rect 450268 3016 465188 579496
rect 465628 3016 480548 579496
rect 480988 3016 495908 579496
rect 496348 3016 511268 579496
rect 511708 3016 526628 579496
rect 527068 3016 541988 579496
rect 542428 3016 557348 579496
rect 557788 3016 572708 579496
rect 573148 3016 579348 579496
rect 2380 578 579348 3016
<< labels >>
rlabel metal3 s 578569 236544 579369 236656 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 441728 582153 441840 582953 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 377664 582153 377776 582953 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 313600 582153 313712 582953 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 249536 582153 249648 582953 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 185472 582153 185584 582953 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121408 582153 121520 582953 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 57344 582153 57456 582953 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 576352 800 576464 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 533344 800 533456 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 490336 800 490448 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 578569 280448 579369 280560 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 447328 800 447440 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 404320 800 404432 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 361312 800 361424 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 318304 800 318416 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 275296 800 275408 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 232288 800 232400 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 189280 800 189392 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 146272 800 146384 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 103264 800 103376 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 578569 324352 579369 324464 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 578569 368256 579369 368368 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 578569 412160 579369 412272 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 578569 456064 579369 456176 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 578569 499968 579369 500080 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 578569 543872 579369 543984 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 569856 582153 569968 582953 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 505792 582153 505904 582953 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 578569 6048 579369 6160 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 578569 379232 579369 379344 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 578569 423136 579369 423248 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 578569 467040 579369 467152 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 578569 510944 579369 511056 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 578569 554848 579369 554960 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 553840 582153 553952 582953 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 489776 582153 489888 582953 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 425712 582153 425824 582953 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 361648 582153 361760 582953 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 297584 582153 297696 582953 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 578569 38976 579369 39088 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 233520 582153 233632 582953 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 169456 582153 169568 582953 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105392 582153 105504 582953 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 41328 582153 41440 582953 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 565600 800 565712 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 522592 800 522704 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 479584 800 479696 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 436576 800 436688 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 393568 800 393680 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 350560 800 350672 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 578569 71904 579369 72016 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 307552 800 307664 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 264544 800 264656 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 221536 800 221648 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 178528 800 178640 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 135520 800 135632 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 92512 800 92624 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 60256 800 60368 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 28000 800 28112 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 578569 104832 579369 104944 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 578569 137760 579369 137872 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 578569 170688 579369 170800 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 578569 203616 579369 203728 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 578569 247520 579369 247632 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 578569 291424 579369 291536 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 578569 335328 579369 335440 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 578569 28000 579369 28112 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 578569 401184 579369 401296 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 578569 445088 579369 445200 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 578569 488992 579369 489104 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 578569 532896 579369 533008 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 578569 576800 579369 576912 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 521808 582153 521920 582953 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 457744 582153 457856 582953 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 393680 582153 393792 582953 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 329616 582153 329728 582953 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 265552 582153 265664 582953 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 578569 60928 579369 61040 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 201488 582153 201600 582953 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137424 582153 137536 582953 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 73360 582153 73472 582953 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 9296 582153 9408 582953 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 544096 800 544208 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 501088 800 501200 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 458080 800 458192 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 415072 800 415184 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 372064 800 372176 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 329056 800 329168 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 578569 93856 579369 93968 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 286048 800 286160 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 243040 800 243152 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 200032 800 200144 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 157024 800 157136 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 114016 800 114128 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 71008 800 71120 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 38752 800 38864 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 6496 800 6608 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 578569 126784 579369 126896 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 578569 159712 579369 159824 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 578569 192640 579369 192752 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 578569 225568 579369 225680 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 578569 269472 579369 269584 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 578569 313376 579369 313488 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 578569 357280 579369 357392 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 578569 17024 579369 17136 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 578569 390208 579369 390320 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 578569 434112 579369 434224 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 578569 478016 579369 478128 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 578569 521920 579369 522032 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 578569 565824 579369 565936 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 537824 582153 537936 582953 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 473760 582153 473872 582953 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 409696 582153 409808 582953 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 345632 582153 345744 582953 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 281568 582153 281680 582953 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 578569 49952 579369 50064 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 217504 582153 217616 582953 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 153440 582153 153552 582953 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89376 582153 89488 582953 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 25312 582153 25424 582953 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 554848 800 554960 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 511840 800 511952 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 468832 800 468944 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 425824 800 425936 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 382816 800 382928 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 339808 800 339920 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 578569 82880 579369 82992 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 296800 800 296912 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 253792 800 253904 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 210784 800 210896 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 167776 800 167888 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 124768 800 124880 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 81760 800 81872 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 49504 800 49616 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 17248 800 17360 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 578569 115808 579369 115920 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 578569 148736 579369 148848 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 578569 181664 579369 181776 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 578569 214592 579369 214704 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 578569 258496 579369 258608 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 578569 302400 579369 302512 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 578569 346304 579369 346416 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 204848 0 204960 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 261968 0 262080 800 6 la_data_in[10]
port 145 nsew signal input
rlabel metal2 s 267680 0 267792 800 6 la_data_in[11]
port 146 nsew signal input
rlabel metal2 s 273392 0 273504 800 6 la_data_in[12]
port 147 nsew signal input
rlabel metal2 s 279104 0 279216 800 6 la_data_in[13]
port 148 nsew signal input
rlabel metal2 s 284816 0 284928 800 6 la_data_in[14]
port 149 nsew signal input
rlabel metal2 s 290528 0 290640 800 6 la_data_in[15]
port 150 nsew signal input
rlabel metal2 s 296240 0 296352 800 6 la_data_in[16]
port 151 nsew signal input
rlabel metal2 s 301952 0 302064 800 6 la_data_in[17]
port 152 nsew signal input
rlabel metal2 s 307664 0 307776 800 6 la_data_in[18]
port 153 nsew signal input
rlabel metal2 s 313376 0 313488 800 6 la_data_in[19]
port 154 nsew signal input
rlabel metal2 s 210560 0 210672 800 6 la_data_in[1]
port 155 nsew signal input
rlabel metal2 s 319088 0 319200 800 6 la_data_in[20]
port 156 nsew signal input
rlabel metal2 s 324800 0 324912 800 6 la_data_in[21]
port 157 nsew signal input
rlabel metal2 s 330512 0 330624 800 6 la_data_in[22]
port 158 nsew signal input
rlabel metal2 s 336224 0 336336 800 6 la_data_in[23]
port 159 nsew signal input
rlabel metal2 s 341936 0 342048 800 6 la_data_in[24]
port 160 nsew signal input
rlabel metal2 s 347648 0 347760 800 6 la_data_in[25]
port 161 nsew signal input
rlabel metal2 s 353360 0 353472 800 6 la_data_in[26]
port 162 nsew signal input
rlabel metal2 s 359072 0 359184 800 6 la_data_in[27]
port 163 nsew signal input
rlabel metal2 s 364784 0 364896 800 6 la_data_in[28]
port 164 nsew signal input
rlabel metal2 s 370496 0 370608 800 6 la_data_in[29]
port 165 nsew signal input
rlabel metal2 s 216272 0 216384 800 6 la_data_in[2]
port 166 nsew signal input
rlabel metal2 s 376208 0 376320 800 6 la_data_in[30]
port 167 nsew signal input
rlabel metal2 s 381920 0 382032 800 6 la_data_in[31]
port 168 nsew signal input
rlabel metal2 s 387632 0 387744 800 6 la_data_in[32]
port 169 nsew signal input
rlabel metal2 s 393344 0 393456 800 6 la_data_in[33]
port 170 nsew signal input
rlabel metal2 s 399056 0 399168 800 6 la_data_in[34]
port 171 nsew signal input
rlabel metal2 s 404768 0 404880 800 6 la_data_in[35]
port 172 nsew signal input
rlabel metal2 s 410480 0 410592 800 6 la_data_in[36]
port 173 nsew signal input
rlabel metal2 s 416192 0 416304 800 6 la_data_in[37]
port 174 nsew signal input
rlabel metal2 s 421904 0 422016 800 6 la_data_in[38]
port 175 nsew signal input
rlabel metal2 s 427616 0 427728 800 6 la_data_in[39]
port 176 nsew signal input
rlabel metal2 s 221984 0 222096 800 6 la_data_in[3]
port 177 nsew signal input
rlabel metal2 s 433328 0 433440 800 6 la_data_in[40]
port 178 nsew signal input
rlabel metal2 s 439040 0 439152 800 6 la_data_in[41]
port 179 nsew signal input
rlabel metal2 s 444752 0 444864 800 6 la_data_in[42]
port 180 nsew signal input
rlabel metal2 s 450464 0 450576 800 6 la_data_in[43]
port 181 nsew signal input
rlabel metal2 s 456176 0 456288 800 6 la_data_in[44]
port 182 nsew signal input
rlabel metal2 s 461888 0 462000 800 6 la_data_in[45]
port 183 nsew signal input
rlabel metal2 s 467600 0 467712 800 6 la_data_in[46]
port 184 nsew signal input
rlabel metal2 s 473312 0 473424 800 6 la_data_in[47]
port 185 nsew signal input
rlabel metal2 s 479024 0 479136 800 6 la_data_in[48]
port 186 nsew signal input
rlabel metal2 s 484736 0 484848 800 6 la_data_in[49]
port 187 nsew signal input
rlabel metal2 s 227696 0 227808 800 6 la_data_in[4]
port 188 nsew signal input
rlabel metal2 s 490448 0 490560 800 6 la_data_in[50]
port 189 nsew signal input
rlabel metal2 s 496160 0 496272 800 6 la_data_in[51]
port 190 nsew signal input
rlabel metal2 s 501872 0 501984 800 6 la_data_in[52]
port 191 nsew signal input
rlabel metal2 s 507584 0 507696 800 6 la_data_in[53]
port 192 nsew signal input
rlabel metal2 s 513296 0 513408 800 6 la_data_in[54]
port 193 nsew signal input
rlabel metal2 s 519008 0 519120 800 6 la_data_in[55]
port 194 nsew signal input
rlabel metal2 s 524720 0 524832 800 6 la_data_in[56]
port 195 nsew signal input
rlabel metal2 s 530432 0 530544 800 6 la_data_in[57]
port 196 nsew signal input
rlabel metal2 s 536144 0 536256 800 6 la_data_in[58]
port 197 nsew signal input
rlabel metal2 s 541856 0 541968 800 6 la_data_in[59]
port 198 nsew signal input
rlabel metal2 s 233408 0 233520 800 6 la_data_in[5]
port 199 nsew signal input
rlabel metal2 s 547568 0 547680 800 6 la_data_in[60]
port 200 nsew signal input
rlabel metal2 s 553280 0 553392 800 6 la_data_in[61]
port 201 nsew signal input
rlabel metal2 s 558992 0 559104 800 6 la_data_in[62]
port 202 nsew signal input
rlabel metal2 s 564704 0 564816 800 6 la_data_in[63]
port 203 nsew signal input
rlabel metal2 s 239120 0 239232 800 6 la_data_in[6]
port 204 nsew signal input
rlabel metal2 s 244832 0 244944 800 6 la_data_in[7]
port 205 nsew signal input
rlabel metal2 s 250544 0 250656 800 6 la_data_in[8]
port 206 nsew signal input
rlabel metal2 s 256256 0 256368 800 6 la_data_in[9]
port 207 nsew signal input
rlabel metal2 s 206752 0 206864 800 6 la_data_out[0]
port 208 nsew signal output
rlabel metal2 s 263872 0 263984 800 6 la_data_out[10]
port 209 nsew signal output
rlabel metal2 s 269584 0 269696 800 6 la_data_out[11]
port 210 nsew signal output
rlabel metal2 s 275296 0 275408 800 6 la_data_out[12]
port 211 nsew signal output
rlabel metal2 s 281008 0 281120 800 6 la_data_out[13]
port 212 nsew signal output
rlabel metal2 s 286720 0 286832 800 6 la_data_out[14]
port 213 nsew signal output
rlabel metal2 s 292432 0 292544 800 6 la_data_out[15]
port 214 nsew signal output
rlabel metal2 s 298144 0 298256 800 6 la_data_out[16]
port 215 nsew signal output
rlabel metal2 s 303856 0 303968 800 6 la_data_out[17]
port 216 nsew signal output
rlabel metal2 s 309568 0 309680 800 6 la_data_out[18]
port 217 nsew signal output
rlabel metal2 s 315280 0 315392 800 6 la_data_out[19]
port 218 nsew signal output
rlabel metal2 s 212464 0 212576 800 6 la_data_out[1]
port 219 nsew signal output
rlabel metal2 s 320992 0 321104 800 6 la_data_out[20]
port 220 nsew signal output
rlabel metal2 s 326704 0 326816 800 6 la_data_out[21]
port 221 nsew signal output
rlabel metal2 s 332416 0 332528 800 6 la_data_out[22]
port 222 nsew signal output
rlabel metal2 s 338128 0 338240 800 6 la_data_out[23]
port 223 nsew signal output
rlabel metal2 s 343840 0 343952 800 6 la_data_out[24]
port 224 nsew signal output
rlabel metal2 s 349552 0 349664 800 6 la_data_out[25]
port 225 nsew signal output
rlabel metal2 s 355264 0 355376 800 6 la_data_out[26]
port 226 nsew signal output
rlabel metal2 s 360976 0 361088 800 6 la_data_out[27]
port 227 nsew signal output
rlabel metal2 s 366688 0 366800 800 6 la_data_out[28]
port 228 nsew signal output
rlabel metal2 s 372400 0 372512 800 6 la_data_out[29]
port 229 nsew signal output
rlabel metal2 s 218176 0 218288 800 6 la_data_out[2]
port 230 nsew signal output
rlabel metal2 s 378112 0 378224 800 6 la_data_out[30]
port 231 nsew signal output
rlabel metal2 s 383824 0 383936 800 6 la_data_out[31]
port 232 nsew signal output
rlabel metal2 s 389536 0 389648 800 6 la_data_out[32]
port 233 nsew signal output
rlabel metal2 s 395248 0 395360 800 6 la_data_out[33]
port 234 nsew signal output
rlabel metal2 s 400960 0 401072 800 6 la_data_out[34]
port 235 nsew signal output
rlabel metal2 s 406672 0 406784 800 6 la_data_out[35]
port 236 nsew signal output
rlabel metal2 s 412384 0 412496 800 6 la_data_out[36]
port 237 nsew signal output
rlabel metal2 s 418096 0 418208 800 6 la_data_out[37]
port 238 nsew signal output
rlabel metal2 s 423808 0 423920 800 6 la_data_out[38]
port 239 nsew signal output
rlabel metal2 s 429520 0 429632 800 6 la_data_out[39]
port 240 nsew signal output
rlabel metal2 s 223888 0 224000 800 6 la_data_out[3]
port 241 nsew signal output
rlabel metal2 s 435232 0 435344 800 6 la_data_out[40]
port 242 nsew signal output
rlabel metal2 s 440944 0 441056 800 6 la_data_out[41]
port 243 nsew signal output
rlabel metal2 s 446656 0 446768 800 6 la_data_out[42]
port 244 nsew signal output
rlabel metal2 s 452368 0 452480 800 6 la_data_out[43]
port 245 nsew signal output
rlabel metal2 s 458080 0 458192 800 6 la_data_out[44]
port 246 nsew signal output
rlabel metal2 s 463792 0 463904 800 6 la_data_out[45]
port 247 nsew signal output
rlabel metal2 s 469504 0 469616 800 6 la_data_out[46]
port 248 nsew signal output
rlabel metal2 s 475216 0 475328 800 6 la_data_out[47]
port 249 nsew signal output
rlabel metal2 s 480928 0 481040 800 6 la_data_out[48]
port 250 nsew signal output
rlabel metal2 s 486640 0 486752 800 6 la_data_out[49]
port 251 nsew signal output
rlabel metal2 s 229600 0 229712 800 6 la_data_out[4]
port 252 nsew signal output
rlabel metal2 s 492352 0 492464 800 6 la_data_out[50]
port 253 nsew signal output
rlabel metal2 s 498064 0 498176 800 6 la_data_out[51]
port 254 nsew signal output
rlabel metal2 s 503776 0 503888 800 6 la_data_out[52]
port 255 nsew signal output
rlabel metal2 s 509488 0 509600 800 6 la_data_out[53]
port 256 nsew signal output
rlabel metal2 s 515200 0 515312 800 6 la_data_out[54]
port 257 nsew signal output
rlabel metal2 s 520912 0 521024 800 6 la_data_out[55]
port 258 nsew signal output
rlabel metal2 s 526624 0 526736 800 6 la_data_out[56]
port 259 nsew signal output
rlabel metal2 s 532336 0 532448 800 6 la_data_out[57]
port 260 nsew signal output
rlabel metal2 s 538048 0 538160 800 6 la_data_out[58]
port 261 nsew signal output
rlabel metal2 s 543760 0 543872 800 6 la_data_out[59]
port 262 nsew signal output
rlabel metal2 s 235312 0 235424 800 6 la_data_out[5]
port 263 nsew signal output
rlabel metal2 s 549472 0 549584 800 6 la_data_out[60]
port 264 nsew signal output
rlabel metal2 s 555184 0 555296 800 6 la_data_out[61]
port 265 nsew signal output
rlabel metal2 s 560896 0 561008 800 6 la_data_out[62]
port 266 nsew signal output
rlabel metal2 s 566608 0 566720 800 6 la_data_out[63]
port 267 nsew signal output
rlabel metal2 s 241024 0 241136 800 6 la_data_out[6]
port 268 nsew signal output
rlabel metal2 s 246736 0 246848 800 6 la_data_out[7]
port 269 nsew signal output
rlabel metal2 s 252448 0 252560 800 6 la_data_out[8]
port 270 nsew signal output
rlabel metal2 s 258160 0 258272 800 6 la_data_out[9]
port 271 nsew signal output
rlabel metal2 s 208656 0 208768 800 6 la_oenb[0]
port 272 nsew signal input
rlabel metal2 s 265776 0 265888 800 6 la_oenb[10]
port 273 nsew signal input
rlabel metal2 s 271488 0 271600 800 6 la_oenb[11]
port 274 nsew signal input
rlabel metal2 s 277200 0 277312 800 6 la_oenb[12]
port 275 nsew signal input
rlabel metal2 s 282912 0 283024 800 6 la_oenb[13]
port 276 nsew signal input
rlabel metal2 s 288624 0 288736 800 6 la_oenb[14]
port 277 nsew signal input
rlabel metal2 s 294336 0 294448 800 6 la_oenb[15]
port 278 nsew signal input
rlabel metal2 s 300048 0 300160 800 6 la_oenb[16]
port 279 nsew signal input
rlabel metal2 s 305760 0 305872 800 6 la_oenb[17]
port 280 nsew signal input
rlabel metal2 s 311472 0 311584 800 6 la_oenb[18]
port 281 nsew signal input
rlabel metal2 s 317184 0 317296 800 6 la_oenb[19]
port 282 nsew signal input
rlabel metal2 s 214368 0 214480 800 6 la_oenb[1]
port 283 nsew signal input
rlabel metal2 s 322896 0 323008 800 6 la_oenb[20]
port 284 nsew signal input
rlabel metal2 s 328608 0 328720 800 6 la_oenb[21]
port 285 nsew signal input
rlabel metal2 s 334320 0 334432 800 6 la_oenb[22]
port 286 nsew signal input
rlabel metal2 s 340032 0 340144 800 6 la_oenb[23]
port 287 nsew signal input
rlabel metal2 s 345744 0 345856 800 6 la_oenb[24]
port 288 nsew signal input
rlabel metal2 s 351456 0 351568 800 6 la_oenb[25]
port 289 nsew signal input
rlabel metal2 s 357168 0 357280 800 6 la_oenb[26]
port 290 nsew signal input
rlabel metal2 s 362880 0 362992 800 6 la_oenb[27]
port 291 nsew signal input
rlabel metal2 s 368592 0 368704 800 6 la_oenb[28]
port 292 nsew signal input
rlabel metal2 s 374304 0 374416 800 6 la_oenb[29]
port 293 nsew signal input
rlabel metal2 s 220080 0 220192 800 6 la_oenb[2]
port 294 nsew signal input
rlabel metal2 s 380016 0 380128 800 6 la_oenb[30]
port 295 nsew signal input
rlabel metal2 s 385728 0 385840 800 6 la_oenb[31]
port 296 nsew signal input
rlabel metal2 s 391440 0 391552 800 6 la_oenb[32]
port 297 nsew signal input
rlabel metal2 s 397152 0 397264 800 6 la_oenb[33]
port 298 nsew signal input
rlabel metal2 s 402864 0 402976 800 6 la_oenb[34]
port 299 nsew signal input
rlabel metal2 s 408576 0 408688 800 6 la_oenb[35]
port 300 nsew signal input
rlabel metal2 s 414288 0 414400 800 6 la_oenb[36]
port 301 nsew signal input
rlabel metal2 s 420000 0 420112 800 6 la_oenb[37]
port 302 nsew signal input
rlabel metal2 s 425712 0 425824 800 6 la_oenb[38]
port 303 nsew signal input
rlabel metal2 s 431424 0 431536 800 6 la_oenb[39]
port 304 nsew signal input
rlabel metal2 s 225792 0 225904 800 6 la_oenb[3]
port 305 nsew signal input
rlabel metal2 s 437136 0 437248 800 6 la_oenb[40]
port 306 nsew signal input
rlabel metal2 s 442848 0 442960 800 6 la_oenb[41]
port 307 nsew signal input
rlabel metal2 s 448560 0 448672 800 6 la_oenb[42]
port 308 nsew signal input
rlabel metal2 s 454272 0 454384 800 6 la_oenb[43]
port 309 nsew signal input
rlabel metal2 s 459984 0 460096 800 6 la_oenb[44]
port 310 nsew signal input
rlabel metal2 s 465696 0 465808 800 6 la_oenb[45]
port 311 nsew signal input
rlabel metal2 s 471408 0 471520 800 6 la_oenb[46]
port 312 nsew signal input
rlabel metal2 s 477120 0 477232 800 6 la_oenb[47]
port 313 nsew signal input
rlabel metal2 s 482832 0 482944 800 6 la_oenb[48]
port 314 nsew signal input
rlabel metal2 s 488544 0 488656 800 6 la_oenb[49]
port 315 nsew signal input
rlabel metal2 s 231504 0 231616 800 6 la_oenb[4]
port 316 nsew signal input
rlabel metal2 s 494256 0 494368 800 6 la_oenb[50]
port 317 nsew signal input
rlabel metal2 s 499968 0 500080 800 6 la_oenb[51]
port 318 nsew signal input
rlabel metal2 s 505680 0 505792 800 6 la_oenb[52]
port 319 nsew signal input
rlabel metal2 s 511392 0 511504 800 6 la_oenb[53]
port 320 nsew signal input
rlabel metal2 s 517104 0 517216 800 6 la_oenb[54]
port 321 nsew signal input
rlabel metal2 s 522816 0 522928 800 6 la_oenb[55]
port 322 nsew signal input
rlabel metal2 s 528528 0 528640 800 6 la_oenb[56]
port 323 nsew signal input
rlabel metal2 s 534240 0 534352 800 6 la_oenb[57]
port 324 nsew signal input
rlabel metal2 s 539952 0 540064 800 6 la_oenb[58]
port 325 nsew signal input
rlabel metal2 s 545664 0 545776 800 6 la_oenb[59]
port 326 nsew signal input
rlabel metal2 s 237216 0 237328 800 6 la_oenb[5]
port 327 nsew signal input
rlabel metal2 s 551376 0 551488 800 6 la_oenb[60]
port 328 nsew signal input
rlabel metal2 s 557088 0 557200 800 6 la_oenb[61]
port 329 nsew signal input
rlabel metal2 s 562800 0 562912 800 6 la_oenb[62]
port 330 nsew signal input
rlabel metal2 s 568512 0 568624 800 6 la_oenb[63]
port 331 nsew signal input
rlabel metal2 s 242928 0 243040 800 6 la_oenb[6]
port 332 nsew signal input
rlabel metal2 s 248640 0 248752 800 6 la_oenb[7]
port 333 nsew signal input
rlabel metal2 s 254352 0 254464 800 6 la_oenb[8]
port 334 nsew signal input
rlabel metal2 s 260064 0 260176 800 6 la_oenb[9]
port 335 nsew signal input
rlabel metal2 s 570416 0 570528 800 6 user_clock2
port 336 nsew signal input
rlabel metal2 s 572320 0 572432 800 6 user_irq[0]
port 337 nsew signal output
rlabel metal2 s 574224 0 574336 800 6 user_irq[1]
port 338 nsew signal output
rlabel metal2 s 576128 0 576240 800 6 user_irq[2]
port 339 nsew signal output
rlabel metal4 s 4448 3076 4768 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 311648 3076 311968 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 342368 3076 342688 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 373088 3076 373408 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 403808 3076 404128 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 434528 3076 434848 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 465248 3076 465568 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 495968 3076 496288 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 526688 3076 527008 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 557408 3076 557728 579436 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 327008 3076 327328 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 357728 3076 358048 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 388448 3076 388768 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 419168 3076 419488 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 449888 3076 450208 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 480608 3076 480928 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 511328 3076 511648 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 542048 3076 542368 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 572768 3076 573088 579436 6 vss
port 341 nsew ground bidirectional
rlabel metal2 s 3024 0 3136 800 6 wb_clk_i
port 342 nsew signal input
rlabel metal2 s 4928 0 5040 800 6 wb_rst_i
port 343 nsew signal input
rlabel metal2 s 6832 0 6944 800 6 wbs_ack_o
port 344 nsew signal output
rlabel metal2 s 14448 0 14560 800 6 wbs_adr_i[0]
port 345 nsew signal input
rlabel metal2 s 79184 0 79296 800 6 wbs_adr_i[10]
port 346 nsew signal input
rlabel metal2 s 84896 0 85008 800 6 wbs_adr_i[11]
port 347 nsew signal input
rlabel metal2 s 90608 0 90720 800 6 wbs_adr_i[12]
port 348 nsew signal input
rlabel metal2 s 96320 0 96432 800 6 wbs_adr_i[13]
port 349 nsew signal input
rlabel metal2 s 102032 0 102144 800 6 wbs_adr_i[14]
port 350 nsew signal input
rlabel metal2 s 107744 0 107856 800 6 wbs_adr_i[15]
port 351 nsew signal input
rlabel metal2 s 113456 0 113568 800 6 wbs_adr_i[16]
port 352 nsew signal input
rlabel metal2 s 119168 0 119280 800 6 wbs_adr_i[17]
port 353 nsew signal input
rlabel metal2 s 124880 0 124992 800 6 wbs_adr_i[18]
port 354 nsew signal input
rlabel metal2 s 130592 0 130704 800 6 wbs_adr_i[19]
port 355 nsew signal input
rlabel metal2 s 22064 0 22176 800 6 wbs_adr_i[1]
port 356 nsew signal input
rlabel metal2 s 136304 0 136416 800 6 wbs_adr_i[20]
port 357 nsew signal input
rlabel metal2 s 142016 0 142128 800 6 wbs_adr_i[21]
port 358 nsew signal input
rlabel metal2 s 147728 0 147840 800 6 wbs_adr_i[22]
port 359 nsew signal input
rlabel metal2 s 153440 0 153552 800 6 wbs_adr_i[23]
port 360 nsew signal input
rlabel metal2 s 159152 0 159264 800 6 wbs_adr_i[24]
port 361 nsew signal input
rlabel metal2 s 164864 0 164976 800 6 wbs_adr_i[25]
port 362 nsew signal input
rlabel metal2 s 170576 0 170688 800 6 wbs_adr_i[26]
port 363 nsew signal input
rlabel metal2 s 176288 0 176400 800 6 wbs_adr_i[27]
port 364 nsew signal input
rlabel metal2 s 182000 0 182112 800 6 wbs_adr_i[28]
port 365 nsew signal input
rlabel metal2 s 187712 0 187824 800 6 wbs_adr_i[29]
port 366 nsew signal input
rlabel metal2 s 29680 0 29792 800 6 wbs_adr_i[2]
port 367 nsew signal input
rlabel metal2 s 193424 0 193536 800 6 wbs_adr_i[30]
port 368 nsew signal input
rlabel metal2 s 199136 0 199248 800 6 wbs_adr_i[31]
port 369 nsew signal input
rlabel metal2 s 37296 0 37408 800 6 wbs_adr_i[3]
port 370 nsew signal input
rlabel metal2 s 44912 0 45024 800 6 wbs_adr_i[4]
port 371 nsew signal input
rlabel metal2 s 50624 0 50736 800 6 wbs_adr_i[5]
port 372 nsew signal input
rlabel metal2 s 56336 0 56448 800 6 wbs_adr_i[6]
port 373 nsew signal input
rlabel metal2 s 62048 0 62160 800 6 wbs_adr_i[7]
port 374 nsew signal input
rlabel metal2 s 67760 0 67872 800 6 wbs_adr_i[8]
port 375 nsew signal input
rlabel metal2 s 73472 0 73584 800 6 wbs_adr_i[9]
port 376 nsew signal input
rlabel metal2 s 8736 0 8848 800 6 wbs_cyc_i
port 377 nsew signal input
rlabel metal2 s 16352 0 16464 800 6 wbs_dat_i[0]
port 378 nsew signal input
rlabel metal2 s 81088 0 81200 800 6 wbs_dat_i[10]
port 379 nsew signal input
rlabel metal2 s 86800 0 86912 800 6 wbs_dat_i[11]
port 380 nsew signal input
rlabel metal2 s 92512 0 92624 800 6 wbs_dat_i[12]
port 381 nsew signal input
rlabel metal2 s 98224 0 98336 800 6 wbs_dat_i[13]
port 382 nsew signal input
rlabel metal2 s 103936 0 104048 800 6 wbs_dat_i[14]
port 383 nsew signal input
rlabel metal2 s 109648 0 109760 800 6 wbs_dat_i[15]
port 384 nsew signal input
rlabel metal2 s 115360 0 115472 800 6 wbs_dat_i[16]
port 385 nsew signal input
rlabel metal2 s 121072 0 121184 800 6 wbs_dat_i[17]
port 386 nsew signal input
rlabel metal2 s 126784 0 126896 800 6 wbs_dat_i[18]
port 387 nsew signal input
rlabel metal2 s 132496 0 132608 800 6 wbs_dat_i[19]
port 388 nsew signal input
rlabel metal2 s 23968 0 24080 800 6 wbs_dat_i[1]
port 389 nsew signal input
rlabel metal2 s 138208 0 138320 800 6 wbs_dat_i[20]
port 390 nsew signal input
rlabel metal2 s 143920 0 144032 800 6 wbs_dat_i[21]
port 391 nsew signal input
rlabel metal2 s 149632 0 149744 800 6 wbs_dat_i[22]
port 392 nsew signal input
rlabel metal2 s 155344 0 155456 800 6 wbs_dat_i[23]
port 393 nsew signal input
rlabel metal2 s 161056 0 161168 800 6 wbs_dat_i[24]
port 394 nsew signal input
rlabel metal2 s 166768 0 166880 800 6 wbs_dat_i[25]
port 395 nsew signal input
rlabel metal2 s 172480 0 172592 800 6 wbs_dat_i[26]
port 396 nsew signal input
rlabel metal2 s 178192 0 178304 800 6 wbs_dat_i[27]
port 397 nsew signal input
rlabel metal2 s 183904 0 184016 800 6 wbs_dat_i[28]
port 398 nsew signal input
rlabel metal2 s 189616 0 189728 800 6 wbs_dat_i[29]
port 399 nsew signal input
rlabel metal2 s 31584 0 31696 800 6 wbs_dat_i[2]
port 400 nsew signal input
rlabel metal2 s 195328 0 195440 800 6 wbs_dat_i[30]
port 401 nsew signal input
rlabel metal2 s 201040 0 201152 800 6 wbs_dat_i[31]
port 402 nsew signal input
rlabel metal2 s 39200 0 39312 800 6 wbs_dat_i[3]
port 403 nsew signal input
rlabel metal2 s 46816 0 46928 800 6 wbs_dat_i[4]
port 404 nsew signal input
rlabel metal2 s 52528 0 52640 800 6 wbs_dat_i[5]
port 405 nsew signal input
rlabel metal2 s 58240 0 58352 800 6 wbs_dat_i[6]
port 406 nsew signal input
rlabel metal2 s 63952 0 64064 800 6 wbs_dat_i[7]
port 407 nsew signal input
rlabel metal2 s 69664 0 69776 800 6 wbs_dat_i[8]
port 408 nsew signal input
rlabel metal2 s 75376 0 75488 800 6 wbs_dat_i[9]
port 409 nsew signal input
rlabel metal2 s 18256 0 18368 800 6 wbs_dat_o[0]
port 410 nsew signal output
rlabel metal2 s 82992 0 83104 800 6 wbs_dat_o[10]
port 411 nsew signal output
rlabel metal2 s 88704 0 88816 800 6 wbs_dat_o[11]
port 412 nsew signal output
rlabel metal2 s 94416 0 94528 800 6 wbs_dat_o[12]
port 413 nsew signal output
rlabel metal2 s 100128 0 100240 800 6 wbs_dat_o[13]
port 414 nsew signal output
rlabel metal2 s 105840 0 105952 800 6 wbs_dat_o[14]
port 415 nsew signal output
rlabel metal2 s 111552 0 111664 800 6 wbs_dat_o[15]
port 416 nsew signal output
rlabel metal2 s 117264 0 117376 800 6 wbs_dat_o[16]
port 417 nsew signal output
rlabel metal2 s 122976 0 123088 800 6 wbs_dat_o[17]
port 418 nsew signal output
rlabel metal2 s 128688 0 128800 800 6 wbs_dat_o[18]
port 419 nsew signal output
rlabel metal2 s 134400 0 134512 800 6 wbs_dat_o[19]
port 420 nsew signal output
rlabel metal2 s 25872 0 25984 800 6 wbs_dat_o[1]
port 421 nsew signal output
rlabel metal2 s 140112 0 140224 800 6 wbs_dat_o[20]
port 422 nsew signal output
rlabel metal2 s 145824 0 145936 800 6 wbs_dat_o[21]
port 423 nsew signal output
rlabel metal2 s 151536 0 151648 800 6 wbs_dat_o[22]
port 424 nsew signal output
rlabel metal2 s 157248 0 157360 800 6 wbs_dat_o[23]
port 425 nsew signal output
rlabel metal2 s 162960 0 163072 800 6 wbs_dat_o[24]
port 426 nsew signal output
rlabel metal2 s 168672 0 168784 800 6 wbs_dat_o[25]
port 427 nsew signal output
rlabel metal2 s 174384 0 174496 800 6 wbs_dat_o[26]
port 428 nsew signal output
rlabel metal2 s 180096 0 180208 800 6 wbs_dat_o[27]
port 429 nsew signal output
rlabel metal2 s 185808 0 185920 800 6 wbs_dat_o[28]
port 430 nsew signal output
rlabel metal2 s 191520 0 191632 800 6 wbs_dat_o[29]
port 431 nsew signal output
rlabel metal2 s 33488 0 33600 800 6 wbs_dat_o[2]
port 432 nsew signal output
rlabel metal2 s 197232 0 197344 800 6 wbs_dat_o[30]
port 433 nsew signal output
rlabel metal2 s 202944 0 203056 800 6 wbs_dat_o[31]
port 434 nsew signal output
rlabel metal2 s 41104 0 41216 800 6 wbs_dat_o[3]
port 435 nsew signal output
rlabel metal2 s 48720 0 48832 800 6 wbs_dat_o[4]
port 436 nsew signal output
rlabel metal2 s 54432 0 54544 800 6 wbs_dat_o[5]
port 437 nsew signal output
rlabel metal2 s 60144 0 60256 800 6 wbs_dat_o[6]
port 438 nsew signal output
rlabel metal2 s 65856 0 65968 800 6 wbs_dat_o[7]
port 439 nsew signal output
rlabel metal2 s 71568 0 71680 800 6 wbs_dat_o[8]
port 440 nsew signal output
rlabel metal2 s 77280 0 77392 800 6 wbs_dat_o[9]
port 441 nsew signal output
rlabel metal2 s 20160 0 20272 800 6 wbs_sel_i[0]
port 442 nsew signal input
rlabel metal2 s 27776 0 27888 800 6 wbs_sel_i[1]
port 443 nsew signal input
rlabel metal2 s 35392 0 35504 800 6 wbs_sel_i[2]
port 444 nsew signal input
rlabel metal2 s 43008 0 43120 800 6 wbs_sel_i[3]
port 445 nsew signal input
rlabel metal2 s 10640 0 10752 800 6 wbs_stb_i
port 446 nsew signal input
rlabel metal2 s 12544 0 12656 800 6 wbs_we_i
port 447 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 579369 582953
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 261724284
string GDS_FILE /mnt/r/work/Rift2Go_2300_GF180_MPW0/openlane/user_proj_example/runs/22_12_04_14_53/results/signoff/rift2Wrap.magic.gds
string GDS_START 574982
<< end >>

