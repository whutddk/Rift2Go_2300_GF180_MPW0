VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rift2Wrap
  CLASS BLOCK ;
  FOREIGN rift2Wrap ;
  ORIGIN 0.000 0.000 ;
  SIZE 2896.845 BY 2914.765 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1182.720 2896.845 1183.280 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2208.640 2910.765 2209.200 2914.765 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1888.320 2910.765 1888.880 2914.765 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1568.000 2910.765 1568.560 2914.765 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1247.680 2910.765 1248.240 2914.765 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 2910.765 927.920 2914.765 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 2910.765 607.600 2914.765 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 2910.765 287.280 2914.765 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2881.760 4.000 2882.320 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2666.720 4.000 2667.280 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2451.680 4.000 2452.240 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1402.240 2896.845 1402.800 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2236.640 4.000 2237.200 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2021.600 4.000 2022.160 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1806.560 4.000 1807.120 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1591.520 4.000 1592.080 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1376.480 4.000 1377.040 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1161.440 4.000 1162.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 946.400 4.000 946.960 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 731.360 4.000 731.920 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 516.320 4.000 516.880 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1621.760 2896.845 1622.320 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1841.280 2896.845 1841.840 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2060.800 2896.845 2061.360 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2280.320 2896.845 2280.880 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2499.840 2896.845 2500.400 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2719.360 2896.845 2719.920 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2849.280 2910.765 2849.840 2914.765 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2528.960 2910.765 2529.520 2914.765 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 30.240 2896.845 30.800 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1896.160 2896.845 1896.720 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2115.680 2896.845 2116.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2335.200 2896.845 2335.760 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2554.720 2896.845 2555.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2774.240 2896.845 2774.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2769.200 2910.765 2769.760 2914.765 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2448.880 2910.765 2449.440 2914.765 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2128.560 2910.765 2129.120 2914.765 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1808.240 2910.765 1808.800 2914.765 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1487.920 2910.765 1488.480 2914.765 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 194.880 2896.845 195.440 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1167.600 2910.765 1168.160 2914.765 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 847.280 2910.765 847.840 2914.765 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 526.960 2910.765 527.520 2914.765 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.640 2910.765 207.200 2914.765 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2828.000 4.000 2828.560 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2612.960 4.000 2613.520 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2397.920 4.000 2398.480 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2182.880 4.000 2183.440 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1967.840 4.000 1968.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1752.800 4.000 1753.360 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 359.520 2896.845 360.080 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1537.760 4.000 1538.320 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1322.720 4.000 1323.280 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1107.680 4.000 1108.240 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 892.640 4.000 893.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 677.600 4.000 678.160 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 462.560 4.000 463.120 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.280 4.000 301.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 524.160 2896.845 524.720 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 688.800 2896.845 689.360 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 853.440 2896.845 854.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1018.080 2896.845 1018.640 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1237.600 2896.845 1238.160 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1457.120 2896.845 1457.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1676.640 2896.845 1677.200 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 140.000 2896.845 140.560 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2005.920 2896.845 2006.480 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2225.440 2896.845 2226.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2444.960 2896.845 2445.520 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2664.480 2896.845 2665.040 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2884.000 2896.845 2884.560 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2609.040 2910.765 2609.600 2914.765 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2288.720 2910.765 2289.280 2914.765 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1968.400 2910.765 1968.960 2914.765 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1648.080 2910.765 1648.640 2914.765 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1327.760 2910.765 1328.320 2914.765 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 304.640 2896.845 305.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1007.440 2910.765 1008.000 2914.765 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.120 2910.765 687.680 2914.765 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.800 2910.765 367.360 2914.765 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.480 2910.765 47.040 2914.765 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2720.480 4.000 2721.040 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2505.440 4.000 2506.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2290.400 4.000 2290.960 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2075.360 4.000 2075.920 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1860.320 4.000 1860.880 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1645.280 4.000 1645.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 469.280 2896.845 469.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1430.240 4.000 1430.800 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1215.200 4.000 1215.760 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1000.160 4.000 1000.720 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 785.120 4.000 785.680 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 570.080 4.000 570.640 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.040 4.000 355.600 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.760 4.000 194.320 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.480 4.000 33.040 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 633.920 2896.845 634.480 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 798.560 2896.845 799.120 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 963.200 2896.845 963.760 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1127.840 2896.845 1128.400 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1347.360 2896.845 1347.920 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1566.880 2896.845 1567.440 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1786.400 2896.845 1786.960 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 85.120 2896.845 85.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1951.040 2896.845 1951.600 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2170.560 2896.845 2171.120 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2390.080 2896.845 2390.640 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2609.600 2896.845 2610.160 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 2829.120 2896.845 2829.680 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2689.120 2910.765 2689.680 2914.765 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2368.800 2910.765 2369.360 2914.765 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2048.480 2910.765 2049.040 2914.765 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1728.160 2910.765 1728.720 2914.765 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1407.840 2910.765 1408.400 2914.765 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 249.760 2896.845 250.320 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1087.520 2910.765 1088.080 2914.765 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 2910.765 767.760 2914.765 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 2910.765 447.440 2914.765 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 2910.765 127.120 2914.765 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2774.240 4.000 2774.800 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2559.200 4.000 2559.760 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2344.160 4.000 2344.720 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2129.120 4.000 2129.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1914.080 4.000 1914.640 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1699.040 4.000 1699.600 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 414.400 2896.845 414.960 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1484.000 4.000 1484.560 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1268.960 4.000 1269.520 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1053.920 4.000 1054.480 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 838.880 4.000 839.440 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 623.840 4.000 624.400 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 247.520 4.000 248.080 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.240 4.000 86.800 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 579.040 2896.845 579.600 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 743.680 2896.845 744.240 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 908.320 2896.845 908.880 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1072.960 2896.845 1073.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1292.480 2896.845 1293.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1512.000 2896.845 1512.560 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2892.845 1731.520 2896.845 1732.080 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1024.240 0.000 1024.800 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1309.840 0.000 1310.400 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1338.400 0.000 1338.960 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1366.960 0.000 1367.520 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1395.520 0.000 1396.080 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1424.080 0.000 1424.640 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1452.640 0.000 1453.200 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1481.200 0.000 1481.760 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1509.760 0.000 1510.320 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1538.320 0.000 1538.880 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1566.880 0.000 1567.440 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1052.800 0.000 1053.360 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1595.440 0.000 1596.000 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1624.000 0.000 1624.560 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1652.560 0.000 1653.120 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1681.120 0.000 1681.680 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1709.680 0.000 1710.240 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1738.240 0.000 1738.800 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1766.800 0.000 1767.360 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1795.360 0.000 1795.920 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1823.920 0.000 1824.480 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1852.480 0.000 1853.040 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1081.360 0.000 1081.920 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1881.040 0.000 1881.600 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1909.600 0.000 1910.160 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1938.160 0.000 1938.720 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1966.720 0.000 1967.280 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1995.280 0.000 1995.840 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2023.840 0.000 2024.400 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2052.400 0.000 2052.960 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2080.960 0.000 2081.520 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2109.520 0.000 2110.080 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2138.080 0.000 2138.640 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1109.920 0.000 1110.480 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2166.640 0.000 2167.200 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2195.200 0.000 2195.760 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2223.760 0.000 2224.320 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2252.320 0.000 2252.880 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2280.880 0.000 2281.440 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2309.440 0.000 2310.000 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2338.000 0.000 2338.560 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2366.560 0.000 2367.120 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2395.120 0.000 2395.680 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2423.680 0.000 2424.240 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1138.480 0.000 1139.040 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2452.240 0.000 2452.800 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2480.800 0.000 2481.360 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2509.360 0.000 2509.920 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2537.920 0.000 2538.480 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2566.480 0.000 2567.040 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2595.040 0.000 2595.600 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2623.600 0.000 2624.160 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2652.160 0.000 2652.720 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2680.720 0.000 2681.280 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2709.280 0.000 2709.840 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1167.040 0.000 1167.600 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2737.840 0.000 2738.400 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2766.400 0.000 2766.960 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2794.960 0.000 2795.520 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2823.520 0.000 2824.080 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1195.600 0.000 1196.160 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1224.160 0.000 1224.720 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1252.720 0.000 1253.280 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1281.280 0.000 1281.840 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1033.760 0.000 1034.320 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1319.360 0.000 1319.920 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1347.920 0.000 1348.480 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1376.480 0.000 1377.040 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1405.040 0.000 1405.600 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1433.600 0.000 1434.160 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1462.160 0.000 1462.720 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1490.720 0.000 1491.280 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1519.280 0.000 1519.840 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1547.840 0.000 1548.400 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1576.400 0.000 1576.960 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1062.320 0.000 1062.880 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1604.960 0.000 1605.520 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1633.520 0.000 1634.080 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1662.080 0.000 1662.640 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1690.640 0.000 1691.200 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1719.200 0.000 1719.760 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1747.760 0.000 1748.320 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1776.320 0.000 1776.880 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1804.880 0.000 1805.440 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1833.440 0.000 1834.000 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1862.000 0.000 1862.560 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1090.880 0.000 1091.440 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1890.560 0.000 1891.120 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1919.120 0.000 1919.680 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1947.680 0.000 1948.240 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1976.240 0.000 1976.800 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2004.800 0.000 2005.360 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2033.360 0.000 2033.920 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2061.920 0.000 2062.480 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2090.480 0.000 2091.040 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2119.040 0.000 2119.600 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2147.600 0.000 2148.160 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1119.440 0.000 1120.000 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2176.160 0.000 2176.720 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2204.720 0.000 2205.280 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2233.280 0.000 2233.840 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2261.840 0.000 2262.400 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2290.400 0.000 2290.960 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2318.960 0.000 2319.520 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2347.520 0.000 2348.080 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2376.080 0.000 2376.640 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2404.640 0.000 2405.200 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2433.200 0.000 2433.760 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1148.000 0.000 1148.560 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2461.760 0.000 2462.320 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2490.320 0.000 2490.880 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2518.880 0.000 2519.440 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2547.440 0.000 2548.000 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2576.000 0.000 2576.560 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2604.560 0.000 2605.120 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2633.120 0.000 2633.680 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2661.680 0.000 2662.240 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2690.240 0.000 2690.800 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2718.800 0.000 2719.360 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1176.560 0.000 1177.120 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2747.360 0.000 2747.920 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2775.920 0.000 2776.480 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2804.480 0.000 2805.040 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2833.040 0.000 2833.600 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1205.120 0.000 1205.680 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1233.680 0.000 1234.240 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1262.240 0.000 1262.800 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1290.800 0.000 1291.360 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1043.280 0.000 1043.840 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1328.880 0.000 1329.440 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1357.440 0.000 1358.000 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1386.000 0.000 1386.560 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1414.560 0.000 1415.120 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1443.120 0.000 1443.680 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1471.680 0.000 1472.240 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1500.240 0.000 1500.800 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1528.800 0.000 1529.360 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1557.360 0.000 1557.920 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1585.920 0.000 1586.480 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 0.000 1072.400 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1614.480 0.000 1615.040 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1643.040 0.000 1643.600 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1671.600 0.000 1672.160 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1700.160 0.000 1700.720 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1728.720 0.000 1729.280 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 0.000 1757.840 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1785.840 0.000 1786.400 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1814.400 0.000 1814.960 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1842.960 0.000 1843.520 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1871.520 0.000 1872.080 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1100.400 0.000 1100.960 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1900.080 0.000 1900.640 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1928.640 0.000 1929.200 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1957.200 0.000 1957.760 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1985.760 0.000 1986.320 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2014.320 0.000 2014.880 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2042.880 0.000 2043.440 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2071.440 0.000 2072.000 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2100.000 0.000 2100.560 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2128.560 0.000 2129.120 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2157.120 0.000 2157.680 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 0.000 1129.520 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2185.680 0.000 2186.240 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2214.240 0.000 2214.800 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2242.800 0.000 2243.360 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2271.360 0.000 2271.920 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2299.920 0.000 2300.480 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2328.480 0.000 2329.040 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2357.040 0.000 2357.600 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2385.600 0.000 2386.160 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2414.160 0.000 2414.720 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2442.720 0.000 2443.280 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1157.520 0.000 1158.080 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2471.280 0.000 2471.840 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2499.840 0.000 2500.400 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2528.400 0.000 2528.960 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2556.960 0.000 2557.520 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2585.520 0.000 2586.080 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2614.080 0.000 2614.640 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2642.640 0.000 2643.200 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2671.200 0.000 2671.760 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2699.760 0.000 2700.320 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2728.320 0.000 2728.880 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 0.000 1186.640 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2756.880 0.000 2757.440 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2785.440 0.000 2786.000 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2814.000 0.000 2814.560 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2842.560 0.000 2843.120 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1214.640 0.000 1215.200 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1243.200 0.000 1243.760 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1271.760 0.000 1272.320 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 0.000 1300.880 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2852.080 0.000 2852.640 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2861.600 0.000 2862.160 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2871.120 0.000 2871.680 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2880.640 0.000 2881.200 4.000 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 2897.180 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 2897.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2863.840 15.380 2865.440 2897.180 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.120 0.000 15.680 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 0.000 25.200 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.160 0.000 34.720 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.240 0.000 72.800 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.920 0.000 396.480 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.040 0.000 453.600 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.160 0.000 510.720 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 0.000 539.280 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.280 0.000 567.840 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 595.840 0.000 596.400 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.400 0.000 624.960 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 652.960 0.000 653.520 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.320 0.000 110.880 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 681.520 0.000 682.080 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 0.000 710.640 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 738.640 0.000 739.200 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 795.760 0.000 796.320 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 0.000 824.880 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 852.880 0.000 853.440 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 0.000 882.000 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.000 0.000 910.560 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 0.000 939.120 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.400 0.000 148.960 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 967.120 0.000 967.680 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 995.680 0.000 996.240 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.480 0.000 187.040 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.560 0.000 225.120 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 0.000 282.240 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 0.000 310.800 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 0.000 339.360 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 0.000 406.000 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.000 0.000 434.560 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 0.000 463.120 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.120 0.000 491.680 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 0.000 520.240 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.240 0.000 548.800 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 576.800 0.000 577.360 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 605.360 0.000 605.920 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 662.480 0.000 663.040 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 691.040 0.000 691.600 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.600 0.000 720.160 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 0.000 748.720 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.720 0.000 777.280 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 805.280 0.000 805.840 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 833.840 0.000 834.400 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.960 0.000 891.520 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 919.520 0.000 920.080 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 948.080 0.000 948.640 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 976.640 0.000 977.200 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1005.200 0.000 1005.760 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.640 0.000 263.200 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 0.000 291.760 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.760 0.000 320.320 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.880 0.000 377.440 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.280 0.000 91.840 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 414.960 0.000 415.520 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 0.000 444.080 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.080 0.000 472.640 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.200 0.000 529.760 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 0.000 558.320 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.320 0.000 586.880 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 643.440 0.000 644.000 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.360 0.000 129.920 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 700.560 0.000 701.120 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 0.000 729.680 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 757.680 0.000 758.240 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 0.000 786.800 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.800 0.000 815.360 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 0.000 843.920 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 871.920 0.000 872.480 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 900.480 0.000 901.040 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 929.040 0.000 929.600 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 0.000 958.160 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.440 0.000 168.000 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 986.160 0.000 986.720 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 0.000 1015.280 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.520 0.000 206.080 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 243.600 0.000 244.160 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.720 0.000 301.280 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.840 0.000 358.400 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 0.000 53.760 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 2895.670 2897.850 ;
      LAYER Metal2 ;
        RECT 4.060 2910.465 46.180 2910.765 ;
        RECT 47.340 2910.465 126.260 2910.765 ;
        RECT 127.420 2910.465 206.340 2910.765 ;
        RECT 207.500 2910.465 286.420 2910.765 ;
        RECT 287.580 2910.465 366.500 2910.765 ;
        RECT 367.660 2910.465 446.580 2910.765 ;
        RECT 447.740 2910.465 526.660 2910.765 ;
        RECT 527.820 2910.465 606.740 2910.765 ;
        RECT 607.900 2910.465 686.820 2910.765 ;
        RECT 687.980 2910.465 766.900 2910.765 ;
        RECT 768.060 2910.465 846.980 2910.765 ;
        RECT 848.140 2910.465 927.060 2910.765 ;
        RECT 928.220 2910.465 1007.140 2910.765 ;
        RECT 1008.300 2910.465 1087.220 2910.765 ;
        RECT 1088.380 2910.465 1167.300 2910.765 ;
        RECT 1168.460 2910.465 1247.380 2910.765 ;
        RECT 1248.540 2910.465 1327.460 2910.765 ;
        RECT 1328.620 2910.465 1407.540 2910.765 ;
        RECT 1408.700 2910.465 1487.620 2910.765 ;
        RECT 1488.780 2910.465 1567.700 2910.765 ;
        RECT 1568.860 2910.465 1647.780 2910.765 ;
        RECT 1648.940 2910.465 1727.860 2910.765 ;
        RECT 1729.020 2910.465 1807.940 2910.765 ;
        RECT 1809.100 2910.465 1888.020 2910.765 ;
        RECT 1889.180 2910.465 1968.100 2910.765 ;
        RECT 1969.260 2910.465 2048.180 2910.765 ;
        RECT 2049.340 2910.465 2128.260 2910.765 ;
        RECT 2129.420 2910.465 2208.340 2910.765 ;
        RECT 2209.500 2910.465 2288.420 2910.765 ;
        RECT 2289.580 2910.465 2368.500 2910.765 ;
        RECT 2369.660 2910.465 2448.580 2910.765 ;
        RECT 2449.740 2910.465 2528.660 2910.765 ;
        RECT 2529.820 2910.465 2608.740 2910.765 ;
        RECT 2609.900 2910.465 2688.820 2910.765 ;
        RECT 2689.980 2910.465 2768.900 2910.765 ;
        RECT 2770.060 2910.465 2848.980 2910.765 ;
        RECT 2850.140 2910.465 2896.740 2910.765 ;
        RECT 4.060 4.300 2896.740 2910.465 ;
        RECT 4.060 1.770 14.820 4.300 ;
        RECT 15.980 1.770 24.340 4.300 ;
        RECT 25.500 1.770 33.860 4.300 ;
        RECT 35.020 1.770 43.380 4.300 ;
        RECT 44.540 1.770 52.900 4.300 ;
        RECT 54.060 1.770 62.420 4.300 ;
        RECT 63.580 1.770 71.940 4.300 ;
        RECT 73.100 1.770 81.460 4.300 ;
        RECT 82.620 1.770 90.980 4.300 ;
        RECT 92.140 1.770 100.500 4.300 ;
        RECT 101.660 1.770 110.020 4.300 ;
        RECT 111.180 1.770 119.540 4.300 ;
        RECT 120.700 1.770 129.060 4.300 ;
        RECT 130.220 1.770 138.580 4.300 ;
        RECT 139.740 1.770 148.100 4.300 ;
        RECT 149.260 1.770 157.620 4.300 ;
        RECT 158.780 1.770 167.140 4.300 ;
        RECT 168.300 1.770 176.660 4.300 ;
        RECT 177.820 1.770 186.180 4.300 ;
        RECT 187.340 1.770 195.700 4.300 ;
        RECT 196.860 1.770 205.220 4.300 ;
        RECT 206.380 1.770 214.740 4.300 ;
        RECT 215.900 1.770 224.260 4.300 ;
        RECT 225.420 1.770 233.780 4.300 ;
        RECT 234.940 1.770 243.300 4.300 ;
        RECT 244.460 1.770 252.820 4.300 ;
        RECT 253.980 1.770 262.340 4.300 ;
        RECT 263.500 1.770 271.860 4.300 ;
        RECT 273.020 1.770 281.380 4.300 ;
        RECT 282.540 1.770 290.900 4.300 ;
        RECT 292.060 1.770 300.420 4.300 ;
        RECT 301.580 1.770 309.940 4.300 ;
        RECT 311.100 1.770 319.460 4.300 ;
        RECT 320.620 1.770 328.980 4.300 ;
        RECT 330.140 1.770 338.500 4.300 ;
        RECT 339.660 1.770 348.020 4.300 ;
        RECT 349.180 1.770 357.540 4.300 ;
        RECT 358.700 1.770 367.060 4.300 ;
        RECT 368.220 1.770 376.580 4.300 ;
        RECT 377.740 1.770 386.100 4.300 ;
        RECT 387.260 1.770 395.620 4.300 ;
        RECT 396.780 1.770 405.140 4.300 ;
        RECT 406.300 1.770 414.660 4.300 ;
        RECT 415.820 1.770 424.180 4.300 ;
        RECT 425.340 1.770 433.700 4.300 ;
        RECT 434.860 1.770 443.220 4.300 ;
        RECT 444.380 1.770 452.740 4.300 ;
        RECT 453.900 1.770 462.260 4.300 ;
        RECT 463.420 1.770 471.780 4.300 ;
        RECT 472.940 1.770 481.300 4.300 ;
        RECT 482.460 1.770 490.820 4.300 ;
        RECT 491.980 1.770 500.340 4.300 ;
        RECT 501.500 1.770 509.860 4.300 ;
        RECT 511.020 1.770 519.380 4.300 ;
        RECT 520.540 1.770 528.900 4.300 ;
        RECT 530.060 1.770 538.420 4.300 ;
        RECT 539.580 1.770 547.940 4.300 ;
        RECT 549.100 1.770 557.460 4.300 ;
        RECT 558.620 1.770 566.980 4.300 ;
        RECT 568.140 1.770 576.500 4.300 ;
        RECT 577.660 1.770 586.020 4.300 ;
        RECT 587.180 1.770 595.540 4.300 ;
        RECT 596.700 1.770 605.060 4.300 ;
        RECT 606.220 1.770 614.580 4.300 ;
        RECT 615.740 1.770 624.100 4.300 ;
        RECT 625.260 1.770 633.620 4.300 ;
        RECT 634.780 1.770 643.140 4.300 ;
        RECT 644.300 1.770 652.660 4.300 ;
        RECT 653.820 1.770 662.180 4.300 ;
        RECT 663.340 1.770 671.700 4.300 ;
        RECT 672.860 1.770 681.220 4.300 ;
        RECT 682.380 1.770 690.740 4.300 ;
        RECT 691.900 1.770 700.260 4.300 ;
        RECT 701.420 1.770 709.780 4.300 ;
        RECT 710.940 1.770 719.300 4.300 ;
        RECT 720.460 1.770 728.820 4.300 ;
        RECT 729.980 1.770 738.340 4.300 ;
        RECT 739.500 1.770 747.860 4.300 ;
        RECT 749.020 1.770 757.380 4.300 ;
        RECT 758.540 1.770 766.900 4.300 ;
        RECT 768.060 1.770 776.420 4.300 ;
        RECT 777.580 1.770 785.940 4.300 ;
        RECT 787.100 1.770 795.460 4.300 ;
        RECT 796.620 1.770 804.980 4.300 ;
        RECT 806.140 1.770 814.500 4.300 ;
        RECT 815.660 1.770 824.020 4.300 ;
        RECT 825.180 1.770 833.540 4.300 ;
        RECT 834.700 1.770 843.060 4.300 ;
        RECT 844.220 1.770 852.580 4.300 ;
        RECT 853.740 1.770 862.100 4.300 ;
        RECT 863.260 1.770 871.620 4.300 ;
        RECT 872.780 1.770 881.140 4.300 ;
        RECT 882.300 1.770 890.660 4.300 ;
        RECT 891.820 1.770 900.180 4.300 ;
        RECT 901.340 1.770 909.700 4.300 ;
        RECT 910.860 1.770 919.220 4.300 ;
        RECT 920.380 1.770 928.740 4.300 ;
        RECT 929.900 1.770 938.260 4.300 ;
        RECT 939.420 1.770 947.780 4.300 ;
        RECT 948.940 1.770 957.300 4.300 ;
        RECT 958.460 1.770 966.820 4.300 ;
        RECT 967.980 1.770 976.340 4.300 ;
        RECT 977.500 1.770 985.860 4.300 ;
        RECT 987.020 1.770 995.380 4.300 ;
        RECT 996.540 1.770 1004.900 4.300 ;
        RECT 1006.060 1.770 1014.420 4.300 ;
        RECT 1015.580 1.770 1023.940 4.300 ;
        RECT 1025.100 1.770 1033.460 4.300 ;
        RECT 1034.620 1.770 1042.980 4.300 ;
        RECT 1044.140 1.770 1052.500 4.300 ;
        RECT 1053.660 1.770 1062.020 4.300 ;
        RECT 1063.180 1.770 1071.540 4.300 ;
        RECT 1072.700 1.770 1081.060 4.300 ;
        RECT 1082.220 1.770 1090.580 4.300 ;
        RECT 1091.740 1.770 1100.100 4.300 ;
        RECT 1101.260 1.770 1109.620 4.300 ;
        RECT 1110.780 1.770 1119.140 4.300 ;
        RECT 1120.300 1.770 1128.660 4.300 ;
        RECT 1129.820 1.770 1138.180 4.300 ;
        RECT 1139.340 1.770 1147.700 4.300 ;
        RECT 1148.860 1.770 1157.220 4.300 ;
        RECT 1158.380 1.770 1166.740 4.300 ;
        RECT 1167.900 1.770 1176.260 4.300 ;
        RECT 1177.420 1.770 1185.780 4.300 ;
        RECT 1186.940 1.770 1195.300 4.300 ;
        RECT 1196.460 1.770 1204.820 4.300 ;
        RECT 1205.980 1.770 1214.340 4.300 ;
        RECT 1215.500 1.770 1223.860 4.300 ;
        RECT 1225.020 1.770 1233.380 4.300 ;
        RECT 1234.540 1.770 1242.900 4.300 ;
        RECT 1244.060 1.770 1252.420 4.300 ;
        RECT 1253.580 1.770 1261.940 4.300 ;
        RECT 1263.100 1.770 1271.460 4.300 ;
        RECT 1272.620 1.770 1280.980 4.300 ;
        RECT 1282.140 1.770 1290.500 4.300 ;
        RECT 1291.660 1.770 1300.020 4.300 ;
        RECT 1301.180 1.770 1309.540 4.300 ;
        RECT 1310.700 1.770 1319.060 4.300 ;
        RECT 1320.220 1.770 1328.580 4.300 ;
        RECT 1329.740 1.770 1338.100 4.300 ;
        RECT 1339.260 1.770 1347.620 4.300 ;
        RECT 1348.780 1.770 1357.140 4.300 ;
        RECT 1358.300 1.770 1366.660 4.300 ;
        RECT 1367.820 1.770 1376.180 4.300 ;
        RECT 1377.340 1.770 1385.700 4.300 ;
        RECT 1386.860 1.770 1395.220 4.300 ;
        RECT 1396.380 1.770 1404.740 4.300 ;
        RECT 1405.900 1.770 1414.260 4.300 ;
        RECT 1415.420 1.770 1423.780 4.300 ;
        RECT 1424.940 1.770 1433.300 4.300 ;
        RECT 1434.460 1.770 1442.820 4.300 ;
        RECT 1443.980 1.770 1452.340 4.300 ;
        RECT 1453.500 1.770 1461.860 4.300 ;
        RECT 1463.020 1.770 1471.380 4.300 ;
        RECT 1472.540 1.770 1480.900 4.300 ;
        RECT 1482.060 1.770 1490.420 4.300 ;
        RECT 1491.580 1.770 1499.940 4.300 ;
        RECT 1501.100 1.770 1509.460 4.300 ;
        RECT 1510.620 1.770 1518.980 4.300 ;
        RECT 1520.140 1.770 1528.500 4.300 ;
        RECT 1529.660 1.770 1538.020 4.300 ;
        RECT 1539.180 1.770 1547.540 4.300 ;
        RECT 1548.700 1.770 1557.060 4.300 ;
        RECT 1558.220 1.770 1566.580 4.300 ;
        RECT 1567.740 1.770 1576.100 4.300 ;
        RECT 1577.260 1.770 1585.620 4.300 ;
        RECT 1586.780 1.770 1595.140 4.300 ;
        RECT 1596.300 1.770 1604.660 4.300 ;
        RECT 1605.820 1.770 1614.180 4.300 ;
        RECT 1615.340 1.770 1623.700 4.300 ;
        RECT 1624.860 1.770 1633.220 4.300 ;
        RECT 1634.380 1.770 1642.740 4.300 ;
        RECT 1643.900 1.770 1652.260 4.300 ;
        RECT 1653.420 1.770 1661.780 4.300 ;
        RECT 1662.940 1.770 1671.300 4.300 ;
        RECT 1672.460 1.770 1680.820 4.300 ;
        RECT 1681.980 1.770 1690.340 4.300 ;
        RECT 1691.500 1.770 1699.860 4.300 ;
        RECT 1701.020 1.770 1709.380 4.300 ;
        RECT 1710.540 1.770 1718.900 4.300 ;
        RECT 1720.060 1.770 1728.420 4.300 ;
        RECT 1729.580 1.770 1737.940 4.300 ;
        RECT 1739.100 1.770 1747.460 4.300 ;
        RECT 1748.620 1.770 1756.980 4.300 ;
        RECT 1758.140 1.770 1766.500 4.300 ;
        RECT 1767.660 1.770 1776.020 4.300 ;
        RECT 1777.180 1.770 1785.540 4.300 ;
        RECT 1786.700 1.770 1795.060 4.300 ;
        RECT 1796.220 1.770 1804.580 4.300 ;
        RECT 1805.740 1.770 1814.100 4.300 ;
        RECT 1815.260 1.770 1823.620 4.300 ;
        RECT 1824.780 1.770 1833.140 4.300 ;
        RECT 1834.300 1.770 1842.660 4.300 ;
        RECT 1843.820 1.770 1852.180 4.300 ;
        RECT 1853.340 1.770 1861.700 4.300 ;
        RECT 1862.860 1.770 1871.220 4.300 ;
        RECT 1872.380 1.770 1880.740 4.300 ;
        RECT 1881.900 1.770 1890.260 4.300 ;
        RECT 1891.420 1.770 1899.780 4.300 ;
        RECT 1900.940 1.770 1909.300 4.300 ;
        RECT 1910.460 1.770 1918.820 4.300 ;
        RECT 1919.980 1.770 1928.340 4.300 ;
        RECT 1929.500 1.770 1937.860 4.300 ;
        RECT 1939.020 1.770 1947.380 4.300 ;
        RECT 1948.540 1.770 1956.900 4.300 ;
        RECT 1958.060 1.770 1966.420 4.300 ;
        RECT 1967.580 1.770 1975.940 4.300 ;
        RECT 1977.100 1.770 1985.460 4.300 ;
        RECT 1986.620 1.770 1994.980 4.300 ;
        RECT 1996.140 1.770 2004.500 4.300 ;
        RECT 2005.660 1.770 2014.020 4.300 ;
        RECT 2015.180 1.770 2023.540 4.300 ;
        RECT 2024.700 1.770 2033.060 4.300 ;
        RECT 2034.220 1.770 2042.580 4.300 ;
        RECT 2043.740 1.770 2052.100 4.300 ;
        RECT 2053.260 1.770 2061.620 4.300 ;
        RECT 2062.780 1.770 2071.140 4.300 ;
        RECT 2072.300 1.770 2080.660 4.300 ;
        RECT 2081.820 1.770 2090.180 4.300 ;
        RECT 2091.340 1.770 2099.700 4.300 ;
        RECT 2100.860 1.770 2109.220 4.300 ;
        RECT 2110.380 1.770 2118.740 4.300 ;
        RECT 2119.900 1.770 2128.260 4.300 ;
        RECT 2129.420 1.770 2137.780 4.300 ;
        RECT 2138.940 1.770 2147.300 4.300 ;
        RECT 2148.460 1.770 2156.820 4.300 ;
        RECT 2157.980 1.770 2166.340 4.300 ;
        RECT 2167.500 1.770 2175.860 4.300 ;
        RECT 2177.020 1.770 2185.380 4.300 ;
        RECT 2186.540 1.770 2194.900 4.300 ;
        RECT 2196.060 1.770 2204.420 4.300 ;
        RECT 2205.580 1.770 2213.940 4.300 ;
        RECT 2215.100 1.770 2223.460 4.300 ;
        RECT 2224.620 1.770 2232.980 4.300 ;
        RECT 2234.140 1.770 2242.500 4.300 ;
        RECT 2243.660 1.770 2252.020 4.300 ;
        RECT 2253.180 1.770 2261.540 4.300 ;
        RECT 2262.700 1.770 2271.060 4.300 ;
        RECT 2272.220 1.770 2280.580 4.300 ;
        RECT 2281.740 1.770 2290.100 4.300 ;
        RECT 2291.260 1.770 2299.620 4.300 ;
        RECT 2300.780 1.770 2309.140 4.300 ;
        RECT 2310.300 1.770 2318.660 4.300 ;
        RECT 2319.820 1.770 2328.180 4.300 ;
        RECT 2329.340 1.770 2337.700 4.300 ;
        RECT 2338.860 1.770 2347.220 4.300 ;
        RECT 2348.380 1.770 2356.740 4.300 ;
        RECT 2357.900 1.770 2366.260 4.300 ;
        RECT 2367.420 1.770 2375.780 4.300 ;
        RECT 2376.940 1.770 2385.300 4.300 ;
        RECT 2386.460 1.770 2394.820 4.300 ;
        RECT 2395.980 1.770 2404.340 4.300 ;
        RECT 2405.500 1.770 2413.860 4.300 ;
        RECT 2415.020 1.770 2423.380 4.300 ;
        RECT 2424.540 1.770 2432.900 4.300 ;
        RECT 2434.060 1.770 2442.420 4.300 ;
        RECT 2443.580 1.770 2451.940 4.300 ;
        RECT 2453.100 1.770 2461.460 4.300 ;
        RECT 2462.620 1.770 2470.980 4.300 ;
        RECT 2472.140 1.770 2480.500 4.300 ;
        RECT 2481.660 1.770 2490.020 4.300 ;
        RECT 2491.180 1.770 2499.540 4.300 ;
        RECT 2500.700 1.770 2509.060 4.300 ;
        RECT 2510.220 1.770 2518.580 4.300 ;
        RECT 2519.740 1.770 2528.100 4.300 ;
        RECT 2529.260 1.770 2537.620 4.300 ;
        RECT 2538.780 1.770 2547.140 4.300 ;
        RECT 2548.300 1.770 2556.660 4.300 ;
        RECT 2557.820 1.770 2566.180 4.300 ;
        RECT 2567.340 1.770 2575.700 4.300 ;
        RECT 2576.860 1.770 2585.220 4.300 ;
        RECT 2586.380 1.770 2594.740 4.300 ;
        RECT 2595.900 1.770 2604.260 4.300 ;
        RECT 2605.420 1.770 2613.780 4.300 ;
        RECT 2614.940 1.770 2623.300 4.300 ;
        RECT 2624.460 1.770 2632.820 4.300 ;
        RECT 2633.980 1.770 2642.340 4.300 ;
        RECT 2643.500 1.770 2651.860 4.300 ;
        RECT 2653.020 1.770 2661.380 4.300 ;
        RECT 2662.540 1.770 2670.900 4.300 ;
        RECT 2672.060 1.770 2680.420 4.300 ;
        RECT 2681.580 1.770 2689.940 4.300 ;
        RECT 2691.100 1.770 2699.460 4.300 ;
        RECT 2700.620 1.770 2708.980 4.300 ;
        RECT 2710.140 1.770 2718.500 4.300 ;
        RECT 2719.660 1.770 2728.020 4.300 ;
        RECT 2729.180 1.770 2737.540 4.300 ;
        RECT 2738.700 1.770 2747.060 4.300 ;
        RECT 2748.220 1.770 2756.580 4.300 ;
        RECT 2757.740 1.770 2766.100 4.300 ;
        RECT 2767.260 1.770 2775.620 4.300 ;
        RECT 2776.780 1.770 2785.140 4.300 ;
        RECT 2786.300 1.770 2794.660 4.300 ;
        RECT 2795.820 1.770 2804.180 4.300 ;
        RECT 2805.340 1.770 2813.700 4.300 ;
        RECT 2814.860 1.770 2823.220 4.300 ;
        RECT 2824.380 1.770 2832.740 4.300 ;
        RECT 2833.900 1.770 2842.260 4.300 ;
        RECT 2843.420 1.770 2851.780 4.300 ;
        RECT 2852.940 1.770 2861.300 4.300 ;
        RECT 2862.460 1.770 2870.820 4.300 ;
        RECT 2871.980 1.770 2880.340 4.300 ;
        RECT 2881.500 1.770 2896.740 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 2884.860 2896.790 2906.260 ;
        RECT 4.000 2883.700 2892.545 2884.860 ;
        RECT 4.000 2882.620 2896.790 2883.700 ;
        RECT 4.300 2881.460 2896.790 2882.620 ;
        RECT 4.000 2829.980 2896.790 2881.460 ;
        RECT 4.000 2828.860 2892.545 2829.980 ;
        RECT 4.300 2828.820 2892.545 2828.860 ;
        RECT 4.300 2827.700 2896.790 2828.820 ;
        RECT 4.000 2775.100 2896.790 2827.700 ;
        RECT 4.300 2773.940 2892.545 2775.100 ;
        RECT 4.000 2721.340 2896.790 2773.940 ;
        RECT 4.300 2720.220 2896.790 2721.340 ;
        RECT 4.300 2720.180 2892.545 2720.220 ;
        RECT 4.000 2719.060 2892.545 2720.180 ;
        RECT 4.000 2667.580 2896.790 2719.060 ;
        RECT 4.300 2666.420 2896.790 2667.580 ;
        RECT 4.000 2665.340 2896.790 2666.420 ;
        RECT 4.000 2664.180 2892.545 2665.340 ;
        RECT 4.000 2613.820 2896.790 2664.180 ;
        RECT 4.300 2612.660 2896.790 2613.820 ;
        RECT 4.000 2610.460 2896.790 2612.660 ;
        RECT 4.000 2609.300 2892.545 2610.460 ;
        RECT 4.000 2560.060 2896.790 2609.300 ;
        RECT 4.300 2558.900 2896.790 2560.060 ;
        RECT 4.000 2555.580 2896.790 2558.900 ;
        RECT 4.000 2554.420 2892.545 2555.580 ;
        RECT 4.000 2506.300 2896.790 2554.420 ;
        RECT 4.300 2505.140 2896.790 2506.300 ;
        RECT 4.000 2500.700 2896.790 2505.140 ;
        RECT 4.000 2499.540 2892.545 2500.700 ;
        RECT 4.000 2452.540 2896.790 2499.540 ;
        RECT 4.300 2451.380 2896.790 2452.540 ;
        RECT 4.000 2445.820 2896.790 2451.380 ;
        RECT 4.000 2444.660 2892.545 2445.820 ;
        RECT 4.000 2398.780 2896.790 2444.660 ;
        RECT 4.300 2397.620 2896.790 2398.780 ;
        RECT 4.000 2390.940 2896.790 2397.620 ;
        RECT 4.000 2389.780 2892.545 2390.940 ;
        RECT 4.000 2345.020 2896.790 2389.780 ;
        RECT 4.300 2343.860 2896.790 2345.020 ;
        RECT 4.000 2336.060 2896.790 2343.860 ;
        RECT 4.000 2334.900 2892.545 2336.060 ;
        RECT 4.000 2291.260 2896.790 2334.900 ;
        RECT 4.300 2290.100 2896.790 2291.260 ;
        RECT 4.000 2281.180 2896.790 2290.100 ;
        RECT 4.000 2280.020 2892.545 2281.180 ;
        RECT 4.000 2237.500 2896.790 2280.020 ;
        RECT 4.300 2236.340 2896.790 2237.500 ;
        RECT 4.000 2226.300 2896.790 2236.340 ;
        RECT 4.000 2225.140 2892.545 2226.300 ;
        RECT 4.000 2183.740 2896.790 2225.140 ;
        RECT 4.300 2182.580 2896.790 2183.740 ;
        RECT 4.000 2171.420 2896.790 2182.580 ;
        RECT 4.000 2170.260 2892.545 2171.420 ;
        RECT 4.000 2129.980 2896.790 2170.260 ;
        RECT 4.300 2128.820 2896.790 2129.980 ;
        RECT 4.000 2116.540 2896.790 2128.820 ;
        RECT 4.000 2115.380 2892.545 2116.540 ;
        RECT 4.000 2076.220 2896.790 2115.380 ;
        RECT 4.300 2075.060 2896.790 2076.220 ;
        RECT 4.000 2061.660 2896.790 2075.060 ;
        RECT 4.000 2060.500 2892.545 2061.660 ;
        RECT 4.000 2022.460 2896.790 2060.500 ;
        RECT 4.300 2021.300 2896.790 2022.460 ;
        RECT 4.000 2006.780 2896.790 2021.300 ;
        RECT 4.000 2005.620 2892.545 2006.780 ;
        RECT 4.000 1968.700 2896.790 2005.620 ;
        RECT 4.300 1967.540 2896.790 1968.700 ;
        RECT 4.000 1951.900 2896.790 1967.540 ;
        RECT 4.000 1950.740 2892.545 1951.900 ;
        RECT 4.000 1914.940 2896.790 1950.740 ;
        RECT 4.300 1913.780 2896.790 1914.940 ;
        RECT 4.000 1897.020 2896.790 1913.780 ;
        RECT 4.000 1895.860 2892.545 1897.020 ;
        RECT 4.000 1861.180 2896.790 1895.860 ;
        RECT 4.300 1860.020 2896.790 1861.180 ;
        RECT 4.000 1842.140 2896.790 1860.020 ;
        RECT 4.000 1840.980 2892.545 1842.140 ;
        RECT 4.000 1807.420 2896.790 1840.980 ;
        RECT 4.300 1806.260 2896.790 1807.420 ;
        RECT 4.000 1787.260 2896.790 1806.260 ;
        RECT 4.000 1786.100 2892.545 1787.260 ;
        RECT 4.000 1753.660 2896.790 1786.100 ;
        RECT 4.300 1752.500 2896.790 1753.660 ;
        RECT 4.000 1732.380 2896.790 1752.500 ;
        RECT 4.000 1731.220 2892.545 1732.380 ;
        RECT 4.000 1699.900 2896.790 1731.220 ;
        RECT 4.300 1698.740 2896.790 1699.900 ;
        RECT 4.000 1677.500 2896.790 1698.740 ;
        RECT 4.000 1676.340 2892.545 1677.500 ;
        RECT 4.000 1646.140 2896.790 1676.340 ;
        RECT 4.300 1644.980 2896.790 1646.140 ;
        RECT 4.000 1622.620 2896.790 1644.980 ;
        RECT 4.000 1621.460 2892.545 1622.620 ;
        RECT 4.000 1592.380 2896.790 1621.460 ;
        RECT 4.300 1591.220 2896.790 1592.380 ;
        RECT 4.000 1567.740 2896.790 1591.220 ;
        RECT 4.000 1566.580 2892.545 1567.740 ;
        RECT 4.000 1538.620 2896.790 1566.580 ;
        RECT 4.300 1537.460 2896.790 1538.620 ;
        RECT 4.000 1512.860 2896.790 1537.460 ;
        RECT 4.000 1511.700 2892.545 1512.860 ;
        RECT 4.000 1484.860 2896.790 1511.700 ;
        RECT 4.300 1483.700 2896.790 1484.860 ;
        RECT 4.000 1457.980 2896.790 1483.700 ;
        RECT 4.000 1456.820 2892.545 1457.980 ;
        RECT 4.000 1431.100 2896.790 1456.820 ;
        RECT 4.300 1429.940 2896.790 1431.100 ;
        RECT 4.000 1403.100 2896.790 1429.940 ;
        RECT 4.000 1401.940 2892.545 1403.100 ;
        RECT 4.000 1377.340 2896.790 1401.940 ;
        RECT 4.300 1376.180 2896.790 1377.340 ;
        RECT 4.000 1348.220 2896.790 1376.180 ;
        RECT 4.000 1347.060 2892.545 1348.220 ;
        RECT 4.000 1323.580 2896.790 1347.060 ;
        RECT 4.300 1322.420 2896.790 1323.580 ;
        RECT 4.000 1293.340 2896.790 1322.420 ;
        RECT 4.000 1292.180 2892.545 1293.340 ;
        RECT 4.000 1269.820 2896.790 1292.180 ;
        RECT 4.300 1268.660 2896.790 1269.820 ;
        RECT 4.000 1238.460 2896.790 1268.660 ;
        RECT 4.000 1237.300 2892.545 1238.460 ;
        RECT 4.000 1216.060 2896.790 1237.300 ;
        RECT 4.300 1214.900 2896.790 1216.060 ;
        RECT 4.000 1183.580 2896.790 1214.900 ;
        RECT 4.000 1182.420 2892.545 1183.580 ;
        RECT 4.000 1162.300 2896.790 1182.420 ;
        RECT 4.300 1161.140 2896.790 1162.300 ;
        RECT 4.000 1128.700 2896.790 1161.140 ;
        RECT 4.000 1127.540 2892.545 1128.700 ;
        RECT 4.000 1108.540 2896.790 1127.540 ;
        RECT 4.300 1107.380 2896.790 1108.540 ;
        RECT 4.000 1073.820 2896.790 1107.380 ;
        RECT 4.000 1072.660 2892.545 1073.820 ;
        RECT 4.000 1054.780 2896.790 1072.660 ;
        RECT 4.300 1053.620 2896.790 1054.780 ;
        RECT 4.000 1018.940 2896.790 1053.620 ;
        RECT 4.000 1017.780 2892.545 1018.940 ;
        RECT 4.000 1001.020 2896.790 1017.780 ;
        RECT 4.300 999.860 2896.790 1001.020 ;
        RECT 4.000 964.060 2896.790 999.860 ;
        RECT 4.000 962.900 2892.545 964.060 ;
        RECT 4.000 947.260 2896.790 962.900 ;
        RECT 4.300 946.100 2896.790 947.260 ;
        RECT 4.000 909.180 2896.790 946.100 ;
        RECT 4.000 908.020 2892.545 909.180 ;
        RECT 4.000 893.500 2896.790 908.020 ;
        RECT 4.300 892.340 2896.790 893.500 ;
        RECT 4.000 854.300 2896.790 892.340 ;
        RECT 4.000 853.140 2892.545 854.300 ;
        RECT 4.000 839.740 2896.790 853.140 ;
        RECT 4.300 838.580 2896.790 839.740 ;
        RECT 4.000 799.420 2896.790 838.580 ;
        RECT 4.000 798.260 2892.545 799.420 ;
        RECT 4.000 785.980 2896.790 798.260 ;
        RECT 4.300 784.820 2896.790 785.980 ;
        RECT 4.000 744.540 2896.790 784.820 ;
        RECT 4.000 743.380 2892.545 744.540 ;
        RECT 4.000 732.220 2896.790 743.380 ;
        RECT 4.300 731.060 2896.790 732.220 ;
        RECT 4.000 689.660 2896.790 731.060 ;
        RECT 4.000 688.500 2892.545 689.660 ;
        RECT 4.000 678.460 2896.790 688.500 ;
        RECT 4.300 677.300 2896.790 678.460 ;
        RECT 4.000 634.780 2896.790 677.300 ;
        RECT 4.000 633.620 2892.545 634.780 ;
        RECT 4.000 624.700 2896.790 633.620 ;
        RECT 4.300 623.540 2896.790 624.700 ;
        RECT 4.000 579.900 2896.790 623.540 ;
        RECT 4.000 578.740 2892.545 579.900 ;
        RECT 4.000 570.940 2896.790 578.740 ;
        RECT 4.300 569.780 2896.790 570.940 ;
        RECT 4.000 525.020 2896.790 569.780 ;
        RECT 4.000 523.860 2892.545 525.020 ;
        RECT 4.000 517.180 2896.790 523.860 ;
        RECT 4.300 516.020 2896.790 517.180 ;
        RECT 4.000 470.140 2896.790 516.020 ;
        RECT 4.000 468.980 2892.545 470.140 ;
        RECT 4.000 463.420 2896.790 468.980 ;
        RECT 4.300 462.260 2896.790 463.420 ;
        RECT 4.000 415.260 2896.790 462.260 ;
        RECT 4.000 414.100 2892.545 415.260 ;
        RECT 4.000 409.660 2896.790 414.100 ;
        RECT 4.300 408.500 2896.790 409.660 ;
        RECT 4.000 360.380 2896.790 408.500 ;
        RECT 4.000 359.220 2892.545 360.380 ;
        RECT 4.000 355.900 2896.790 359.220 ;
        RECT 4.300 354.740 2896.790 355.900 ;
        RECT 4.000 305.500 2896.790 354.740 ;
        RECT 4.000 304.340 2892.545 305.500 ;
        RECT 4.000 302.140 2896.790 304.340 ;
        RECT 4.300 300.980 2896.790 302.140 ;
        RECT 4.000 250.620 2896.790 300.980 ;
        RECT 4.000 249.460 2892.545 250.620 ;
        RECT 4.000 248.380 2896.790 249.460 ;
        RECT 4.300 247.220 2896.790 248.380 ;
        RECT 4.000 195.740 2896.790 247.220 ;
        RECT 4.000 194.620 2892.545 195.740 ;
        RECT 4.300 194.580 2892.545 194.620 ;
        RECT 4.300 193.460 2896.790 194.580 ;
        RECT 4.000 140.860 2896.790 193.460 ;
        RECT 4.300 139.700 2892.545 140.860 ;
        RECT 4.000 87.100 2896.790 139.700 ;
        RECT 4.300 85.980 2896.790 87.100 ;
        RECT 4.300 85.940 2892.545 85.980 ;
        RECT 4.000 84.820 2892.545 85.940 ;
        RECT 4.000 33.340 2896.790 84.820 ;
        RECT 4.300 32.180 2896.790 33.340 ;
        RECT 4.000 31.100 2896.790 32.180 ;
        RECT 4.000 29.940 2892.545 31.100 ;
        RECT 4.000 1.820 2896.790 29.940 ;
      LAYER Metal4 ;
        RECT 11.900 2897.480 2896.740 2905.750 ;
        RECT 11.900 15.080 21.940 2897.480 ;
        RECT 24.140 15.080 98.740 2897.480 ;
        RECT 100.940 15.080 175.540 2897.480 ;
        RECT 177.740 15.080 252.340 2897.480 ;
        RECT 254.540 15.080 329.140 2897.480 ;
        RECT 331.340 15.080 405.940 2897.480 ;
        RECT 408.140 15.080 482.740 2897.480 ;
        RECT 484.940 15.080 559.540 2897.480 ;
        RECT 561.740 15.080 636.340 2897.480 ;
        RECT 638.540 15.080 713.140 2897.480 ;
        RECT 715.340 15.080 789.940 2897.480 ;
        RECT 792.140 15.080 866.740 2897.480 ;
        RECT 868.940 15.080 943.540 2897.480 ;
        RECT 945.740 15.080 1020.340 2897.480 ;
        RECT 1022.540 15.080 1097.140 2897.480 ;
        RECT 1099.340 15.080 1173.940 2897.480 ;
        RECT 1176.140 15.080 1250.740 2897.480 ;
        RECT 1252.940 15.080 1327.540 2897.480 ;
        RECT 1329.740 15.080 1404.340 2897.480 ;
        RECT 1406.540 15.080 1481.140 2897.480 ;
        RECT 1483.340 15.080 1557.940 2897.480 ;
        RECT 1560.140 15.080 1634.740 2897.480 ;
        RECT 1636.940 15.080 1711.540 2897.480 ;
        RECT 1713.740 15.080 1788.340 2897.480 ;
        RECT 1790.540 15.080 1865.140 2897.480 ;
        RECT 1867.340 15.080 1941.940 2897.480 ;
        RECT 1944.140 15.080 2018.740 2897.480 ;
        RECT 2020.940 15.080 2095.540 2897.480 ;
        RECT 2097.740 15.080 2172.340 2897.480 ;
        RECT 2174.540 15.080 2249.140 2897.480 ;
        RECT 2251.340 15.080 2325.940 2897.480 ;
        RECT 2328.140 15.080 2402.740 2897.480 ;
        RECT 2404.940 15.080 2479.540 2897.480 ;
        RECT 2481.740 15.080 2556.340 2897.480 ;
        RECT 2558.540 15.080 2633.140 2897.480 ;
        RECT 2635.340 15.080 2709.940 2897.480 ;
        RECT 2712.140 15.080 2786.740 2897.480 ;
        RECT 2788.940 15.080 2863.540 2897.480 ;
        RECT 2865.740 15.080 2896.740 2897.480 ;
        RECT 11.900 2.890 2896.740 15.080 ;
  END
END rift2Wrap
END LIBRARY

